�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?PbM���X   coef0q	G        X   tolq
G?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�C�9�n��?xL�S@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?PbM���X   support_q3hhK �q4h�q5Rq6(KM
�q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B(           	                                 '   -   /   0   3   5   6   :   @   A   B   D   F   G   L   M   O   P   S   T   U   W   X   Y   Z   `   c   e   h   m   n   o   p   r   u   w   x   y   {   |   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �               
                     !  #  )  *  ,  /  1  2  4  5  8  <  >  B  G  H  K  T  Z  ]  _  b  d  e  f  g  h  i  k  l  m  n  o  p  q  r  u  v  w  x  y  }    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �             	  
                !   %   C   V   j   q   s   �   �   �   �   �   �   �   �   �   �       0  7  A  F  I  S  �  �  �  �  �  �  �  �  �      q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KM
K�qBh"�B�)  s����`�?�0�0�?��e�s��?���]�(�?�������?0.Ba��?.�袋.@�
�l�?haz�g�?      �?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?T�.�n��?�-�׮�?H{����?������?P���Q�?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?F}�p �?������?N6����?\����?ffffff�?��ԩ/��?AR˔���?JL �F�?�>,��?�������?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?"K�_y�?���,d�?���<�?jhɬ�?�Q���?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?lv��?*.�u��?m�����?O�<�"�?!��Q��?-����?ӟ���?���;<�?�׷0���?�Q����?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?L�|9��?m���X��?�B�q��?����:.�?833333�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?e�F-��?�������?���:%�?V���g�?ףp=
�?@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?,"�j�%�?,-----�?'狗�8�?�`�����?133333�?U@�'��?�x+�R�??dM2_�?�(S�\��?�(\�����8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?/9(��?.�袋.
@�*����?�������?�������?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?濸����?r���0�?,�C ^��?5���4�?���(\��?톘��=�?+P�W
��?���gk�?�������?Z���(\�?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�ۇA�?��*�3��?���R�]�?AA�?��(\���?�п�cX�?���؜��?��{�z��?�F��?_fffff�?��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�??V�)��?_�_��?      �?��B�
�?�G�z�?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��2���?���?��</�b�?�ռY͛�?H�z�G�?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?���?�m۶m�@��X)�O�?�\.�?)\���(�?���e��?I��/�?i�(�U�?�VC��?T���Q�?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?R8�u�?S{���?��,�1�?:�oO�$�? �G�z������?1bĈ�?��6-f�?�Ab�k�?�������?�>����?      �?0`z��Q�?'u_�?�p=
ף�?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff���,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?�u����?�wK�?��?�ef���?tT����?�z�G��?
��\���?��\AL��?)us�?      �?433333�?���g
�?&���^B@���X^�?��FS���?G�z�G�?�h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?�qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?(� .b��?�k�S��?��F����?���w���? �G�z�?fo/���?/����?'N`�4��?��3���?�������s��&�?(W�7�?���xW�?B�HV��?��(\���?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�2�j���?     �?u�;�F�?�$I�$I�?�z�G��?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�
>U�?
ŭP�
�?Pf�i���? i]���?�G�z��?:+��?NB�3�?Ci!��?r�q��?Y���(\�?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?��p����?      �?��e�N�?�������?R���Q@�4����?�%����?�J:��?v{�e��?���(\��?��bK��?�/��/��?T��cP��?.Ԝ��?�Q����?��9���?�e���?��G��\�?�����\�?���(\��?8����?�gS��=�?�~��H�?�Vi�_�?�������?@i���?P��O���?�k�9���?��U�^�?(\���(�?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?aC�����?     �?J�.����?"1ogH��?��(\���?Ե7�rL�?�l��l��?���'��?��E���?��G�z���מ���?�i�i�?Q�XW��?�R�~���?      �?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?g�\���?�����?��񍔎�?����.��?�G�z�?�}��?       @j��_�?��¯�D�?�(\����?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿Un����?�������?#�R���?]�����?�Q�����%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�C����?�������?A�ra���?�@۽U��?���Q��?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?�X$����?L�:,��?&����?G�N��?\���(�?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?��h�D��?��P��9�?�1$0��?}��O���?833333�?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?��״��?Ѻ���@��O��?����T�?���(\��?��j�G�?u�5�o��?���d��?�~��?�G�z��?:N�1��?G�:y�?Y<�&!�?F����?��(\���?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?������?������?�X^o�?��<t/�?H�z�G�?4s���?�����?/z�V�4�?~"����?H�z�G�?+e��R�?pА����?�_P�
�?���譺�?��(\����܎h�?��/�$�?�p\��?���6�?���(\��?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?ϙΔ�?a#@i��?M��d�?��,��?      �?evoƃ��?�q�u�?�)���R�?t������?0\���(�?L�Q���?����S��? 0 ��?4և����?433333�?_i�"�?VUUUU��?��i��?)\���(�?�������?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=���t�j�?��qg	��?d���1�?(�)��;�?�������?�T����?Z7�"�u@m�����?����T�?�������?�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�W���?{�n��?	sG�h��?в�9��?��(\���?[��`��?ك2�*j�?� �;��?�������?�(\����?��I��?      �?	)�L��?ڟ�!T�?��G�z���0k��(�?�Iݗ�V�?���Y&�?���?�?      �?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿?d~-��?�u�����?����2�?� ?7��?      �?E�X9�x�?-��,�?)=��'�?��0���?�Q����?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?�O�<�?������@uq_�E�?��$2��?H�z�G�?�83���?�{Nm{�?�F�� �?�������?P���Q�?3�J���?�F�tj�?^���i��?�
� ��?�Q����?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?O�TE���?�(፦@��x�b�?��RJ)��?�������?f��UJ��?�!XG��?�����?����vW�?8
ףp=��[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�_����?      @����,��?[�o�W��?���Q��?8P��A��?�\;0��?<b���e�?y{�X�?      �?I��q��?�'iq��?�&��?#�����?�Q����?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?0	�`���?o�vu�?N�� V�?��X���?��Q���?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?mӞ��?#��~j��?�1?��l�?��i���?�Q����?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?�h�(���?����?�3��=�?g�=���?�������?��zZ �?&jW�v%�?t���?X`��?!��Q��?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?�d����?���-���?_l�9��?L��N���?P���Q�?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�?;�H�r��?W�rCH�?��A�^�?�����?(\���(�?�G,���?�	����?���R{�?��?�c��?���Q��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��aJ��?��˝��?�D�y�?�$���?���(\� @u�-BK�?��T��K�?��x���?>���~��?���Q��?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?:����?�5��P�?v$����?;�;��?أp=
��?��]��S�?�z�����?����?1�0��?(\���(�?9gήc��?�Z$�R��?������?�/��/��?033333�6%�M���?���s @N�|ҍV�?e�e��?�������? ��2�?S�n0�?���&�_�?I%�e��?�������?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?�m�02��?;r����?���	���?����<�?��(\���?�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?|A� *��?�袋.�@��k{�?W�+���?H�z�G�?��X��?�Kh/��?�f i5�?*g���?���Q��?���X �?�\�\�?6#�|a�?>6:8���?P���Q�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp�X���A�?������ @<�z^��?C���,�?�������?��{G�?����S�?Y�_��?�����B�?֣p=
��?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�!ފ�?c����?��J%%�?��(\���?�G�z�?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?əPB�?��.���?gL0�h�?l��(�?ףp=
�?�n��?�3_�g��?����B�?`V�4[s�?`fffff����/����?���T4�?h�v�Q�?�����? ףp=
���L���z�?X�O���?��F�{�?!���c��?�(\����?��m��?����?&z`�5�?2u�=�S�?      �?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?
��Y0�?�G*;�?      �?������?��Q��?/������?�k��%�?���g���?8S����?�G�z���0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?~�aE�?"�z\��?�R����?I��/�?.\���(�?`���`��?���-��?����w�?��-�jL�?��(\��ſ�X��S��?      �?Ѹ�U�?1�0��?���Q���r>bܘ�?��MmjS�?e�����?|1����?���(\��?��B\&�?�n0E>��?���L�?2 K��?�(\����?q�ک��?      @���<X�?��=���?333333�?����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?P@��}�?��k���?      �?�J���?�������?F��W~�?��f=Q��?�����?DDDDDD�?P���Q�?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?����g��?�]����?P�øW�?v�=H]��?��Q���?auȒ���?�v%jW�@��s5��?`����?�Q����?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?����?���a���?Û�P�?�`8wC�?P���Q�?l,����?gH���?���2G�?v�A����?�z�G��?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?����?��R�y�?�����?�s@ڦ�?�p=
ף�?������?�~H���?U��oW�?��S�r
�?
ףp=
�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?D���Oz�?PuPu�?      �?٫��J�?���Q��?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?*�fV=�?'���?<��v��?ZLg1���?�������?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?����8��?��*H�?>���h�?�؊���?$\���(�?�����?)�����?�s�H�?�u�y��?�G�z�?����-�?��L��L@;K�*�O�?��
��?�������?�wF�?��D'�?6������?�_�_�?�������?�������?�m����?G��|���?E4Z����?�z�G��?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?���6���?�w���?zkfkl��?�k(���?      @tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�ݭ����?yþ�\�?�CM`��?�w��K�?�p=
��?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?�'���?�*H^�?�����?Oozӛ��?,\���(�?�S�����?���NV��?��=��?^���?��Q�@@�X兞�?f���?����15�?�>��?��Q���?P��-��?�NV�#�?8��m���?�;�#�?333333@�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?5~�lk��?u32"��?8����j�?�����?�z�G��?�q� .�?��"E��?�V���2�?�^�^�?�G�z�?��]���?[�[�@�{�q�?.q����?���Q��?��1���?wF]�K��?={��?������?�Q����?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?ӏK�K�?��{���?���S��?{���g�?P���Q�?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?�p�|���?���)��?^�3���?h�J� :�?�Q����?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?qCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�   (   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM
�qPh"�BP  歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��dS����{�歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��d�~���I�歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��
0gu�H�歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M��歏�M�����8+��@���8+��@���8+��@�>���@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@h	�%c��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@UZ����w@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@���8+��@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�C��_��$@qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�CQ\E����q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�C?`��s��qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�C��_��$�qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM
�qvh"�BP  歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@dS����{@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@d�~���I@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@
0gu�H@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@歏�M�@���8+������8+������8+����>�������8+������8+������8+������8+������8+������8+������8+���h	�%c������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+���UZ����w����8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+������8+���qwtqxbX   _sklearn_versionqyX   0.21.3qzub.