�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?6��C-X   coef0q	G        X   tolq
G?PbM���X   CqKX   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�C?P����?'M�4i�@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?6��C-X   support_q3hhK �q4h�q5Rq6(KM�q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B8                           	   
                                                                !   "   #   $   %   &   '   (   )   +   ,   .   0   1   2   3   4   5   7   9   ;   <   >   ?   A   B   C   D   E   F   G   H   I   J   K   L   M   N   O   P   Q   R   S   T   U   Z   [   \   ]   ^   _   `   a   b   c   d   e   f   g   h   i   j   k   n   o   p   s   t   u   v   w   x   y   z   {   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                  	  
                                             !  "  #  $  %  &  '  (  *  +  -  .  0  1  2  3  4  5  6  7  8  9  :  ;  <  =  >  ?  @  B  C  E  F  G  H  I  J  K  L  M  N  O  P  Q  R  T  U  V  W  Y  Z  [  \  ^  _  `  a  b  c  f  g  h  i  j  k  l  m  n  p  q  r  s  t  u  w  x  y  z  {  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                     	  
                 *   -   /   6   8   :   =   @   V   W   X   Y   l   m   q   r   |   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �         )  ,  /  A  D  S  X  ]  d  e  o  v  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KMK�qBh"�B0R  ���ʦ�?�6f�@��?�~�ϓ�?FM0��>�?�G�z�@F_L�D��?:��8���?�\�]�G�?l�����?������ @s����`�?�0�0�?��e�s��?���]�(�?�������?�&>�K��?��D/ڷ�?$�A��?�8����?֣p=
�@Eb���?��Y@�H�?�|��X.�?�������?��Q��	@��=�9�?�[��"e�?�+U��R�?�Gq�>�?��Q���?0.Ba��?.�袋.@�
�l�?haz�g�?      �?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?T�.�n��?�-�׮�?H{����?������?P���Q�?�jǊ��?������?<�7b��?"�r����?أp=
�	@��H��?�z�G�?G��ֳ�?
݋н�?R���Q@�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?F}�p �?������?N6����?\����?ffffff�?*�fV=�?'���?<��v��?ZLg1���?�������?��ԩ/��?AR˔���?JL �F�?�>,��?�������?E��.��?5�\�`��?���nD�?P��n��?�(\���@�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?������?�{�D!�?�l.�VP�?�2��h.�?)\���(@���*�_�?۶m۶m�?E������?�n���?�p=
ף@0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?"K�_y�?���,d�?���<�?jhɬ�?�Q���?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?9�KO���? ���?R-ŭX�?X�,)D�?\���(\@�!K���?)^ ���?u�`6�?���j��?q=
ףp�?^���*�?Z5�Uc[�?���l��?Ҏ#��?�Q���?R�p,C.�?������?��U�	��?n��x�>�?��Q��@�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?����?��Pp%��?kub�Q�?̟�Ѐ%�?������񿖨��8��?��*H�?>���h�?�؊���?$\���(�?���#�?})�Z�?d#D:��?��;�?��(\��	@Sle�%�?Q��h��?j鱊 ��?��(C��?efffff@�Fm�}�?�/Rm���?q�Q>	�?ݫ`���?=
ףp=@�����?)�����?�s�H�?�u�y��?�G�z�?w��{���?)�b���?z9��E�?�0��=)�?�������-����?ӟ���?���;<�?�׷0���?�Q����?Qn�p&�?�؉�؉�?�*����?��M�`�?�p=
ף@������?S"�?e8����?�^�6���?�p=
ף@�r*��?z�Ha��?��R����?�{mĺ��?���Q�濔y]>d�?g;>)7�?�Ǭ�NR�?&H-/|�?=
ףp=
@i�+s�?333333�?`�>��R�?��.���?q=
ףp@Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@Q�ps[-�?#N�	���?�[�����?��)��
�?������@e�F-��?�������?���:%�?V���g�?ףp=
�?EÓ���?�����?�&z��V�?WUUUU��?���(\�@@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?�t&����?��(��(�?�^mSz��?g�Bg�B�?������@�Dz�:�?�=��!�?���f�?�%��}'�?�p=
ף@x����v�?4H�4H��?�)~�r��?���Kh�?�p=
ףпm�<�?     �?�������?A�zy3A�?{�G�z
@���,��?ى�؉��?��� W��?{�G�z�?*\���(@���E�]�?WUUUUU�?��o3��?p-ܴ�?��Q��@U@�'��?�x+�R�??dM2_�?�(S�\��?�(\�����8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?����-�?��L��L@;K�*�O�?��
��?�������?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?�����?IM0��>�?��I��?�h�k��? R���ѿ/9(��?.�袋.
@�*����?�������?�������?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?��}��?	�#Q�?F�c[�~�?A�V�{�?��Q��@Se�;f�?h����@A�j�}��?�WJ�B��?S���Q @��Zb��?��+x���?� �Y]��?����?hfffff@��;�l�?��{����?��`|��?���!�?@\���(̿濸����?r���0�?,�C ^��?5���4�?���(\��?톘��=�?+P�W
��?���gk�?�������?Z���(\�?��y����?I`�:�?�5G��`�?4h��J�?      п�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�ۇA�?��*�3��?���R�]�?AA�?��(\���?Um�����?�t��N��?�;1��?_�1yo|�?r=
ףp@�@��+W�?��)o���?�߾���?      �?������@�п�cX�?���؜��?��{�z��?�F��?_fffff�?��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�??V�)��?_�_��?      �?��B�
�?�G�z�?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?���Y�?�	g�	g�?ya��w�?!s��2�?�p=
ף@r6]����?�������?�	��6f�?���3$��?H�z�G@oCӱ�>�?Y�eY�e�?�}{�:��?�p'�p'�?������@S\�C{��?5�rO#,�?64�����?�|�G�j�?ףp=
�@<�	��-�?�U'�*6�?4�(�e�?�>���?֣p=
�	@��2���?���?��</�b�?�ռY͛�?H�z�G�?¶�F�s�?0w�fs�?)���k�?y�!���?{�G�z@48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?��sr��?��3���?�V��?��~5&�? ףp=
׿���?�m۶m�@��X)�O�?�\.�?)\���(�?dwl���?d�fI�m�?��W�6\�?=]�:��?)\���(
@\�����?�3�u�?�d�yv6�?f����?���(\�ҿ���e��?I��/�?i�(�U�?�VC��?T���Q�?�4��
:�?(6$�)G�?(��J+z�?v��4��?���(\�@�������?�m����?G��|���?E4Z����?�z�G��?W['s�,�?E�JԮD�?��K�y�?��J�[��?r=
ףp@R8�u�?S{���?��,�1�?:�oO�$�? �G�z������?1bĈ�?��6-f�?�Ab�k�?�������?�>����?      �?0`z��Q�?'u_�?�p=
ף�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?C�Z����?�Nu�w��?��سX��?�R:CW��?H�z�G@�u����?�wK�?��?�ef���?tT����?�z�G��?
��\���?��\AL��?)us�?      �?433333�?���g
�?&���^B@���X^�?��FS���?G�z�G�?��S��?I�$I�$�?�����?���w��?�������?�h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?�4~���?h}�}-�?	+��]��?�ܽ*���?�Q���	@�$�vQ�?����?dȇ���?�?2�խ�?*\���(@����?;�;��?�(N��?�	F��?������@���� �?�$I�$I@W�G#��?"1ogH��?ffffff�?�qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?O@���?ffffff�??w��a�?�A���?��Q���?���J�&�?J)��RJ�?lj�I�#�?�Y�6���?�(\���
@�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?r�2�F�?�zۜ��?z!I�,�?c[:��c�?�p=
ף@M%����?�:�ֆi�??��!i�?��8��8�?���Q��?�'��|-�?HT�n��?^����,�?#e�����?�(\���
@(� .b��?�k�S��?��F����?���w���? �G�z�?
��@��?���Қ�?'::V�e�?��JR�?������	@�Ĭ~��?��Q���?>s=��^�?�����?�(\����?fo/���?/����?'N`�4��?��3���?�������:�X{��?���.{�?P�l�V��?'��,�?      @s��&�?(W�7�?���xW�?B�HV��?��(\���?}��Yc��?���_��?+��6rl�?W�m���?�G�z�	@�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�2�j���?     �?u�;�F�?�$I�$I�?�z�G��?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?b�+d�&�?�L�w�?U�&xl�?=��k�?�(\���
@����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?�
>U�?
ŭP�
�?Pf�i���? i]���?�G�z��?C�oB��?      �??��(b-�?b�1`�?433333@9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?��p����?      �?��e�N�?�������?R���Q@��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?G��?�����?�8�҂�?K0�|w�?
ףp=
@K�^�/�?(✭��?.�, �y�?!z|��?R���Q@*�zHb�?xwwwww�?Ў���J�?캮뺮�?\���(\@�Ni�3�?�l�����?��+���?�S�n�?!��Q��?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?�\7z�?���"��?����}�?7�j�?H�z�G@��bK��?�/��/��?T��cP��?.Ԝ��?�Q����?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?��9���?�e���?��G��\�?�����\�?���(\��?�ꍑ��?�h�����?Xn�e�w�?��:X���?�G�z�@8����?�gS��=�?�~��H�?�Vi�_�?�������?��(��?7�Y�"�?ޤ�=%�?{�!���?���Q� @@i���?P��O���?�k�9���?��U�^�?(\���(�?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?aC�����?     �?J�.����?"1ogH��?��(\���?Ե7�rL�?�l��l��?���'��?��E���?��G�z��(1B���?b'vb'v�?s�ӭ��? �R{���?H�z�G@g�\���?�����?��񍔎�?����.��?�G�z�?��_O�?��G��=�?�!|����?L��7���?033333@)��h��?UUUUUU�?�����g�?�X>b��?���Q��?� �9�$�?h���Q��?�3�s�?�B#�E�?��Q�@�}��?       @j��_�?��¯�D�?�(\����?�$�l���?d!Y�B�?k���?"�?d�*|��? ףp=
׿ 3`���?���P��?�D�e'~�?�]���?{�G�z@9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?�p^��m�?tT����? ����?����x�?���(\�
@��;4��?WUUUUU�?��J�l�?W�m���?H�z�G@���6���?�w���?zkfkl��?�k(���?      @�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿'�CU$
�?      �?�t�U�%�?.�#EC�?��Q�@Un����?�������?#�R���?]�����?�Q�����%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�C����?�������?A�ra���?�@۽U��?���Q��?�y�]��?]�)~I��?��@��[�?�{����?���(\�@���~�?9"�P9�?<O�����?!������?���(\��?:M�]��?HA@s}�?g0�d��?��7���?\���(\@1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?�X$����?L�:,��?&����?G�N��?\���(�?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@�x�\�?��2����?ؔ�
&w�?      �?أp=
�@�D̥�
�?�Zk����?��iz�?���\��?��Q���?I)i���?�{0�I��?KU���?�X�����?@
ףp=�e�@���?�E�=?2�?Pr^u���?O!�i��?ףp=
�@-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?�i����?T����|�?�;x�]z�?,d!Y��?P���Q�?��L��?�q�q�?G`3�!�?O���t:�?R���Q@��h�D��?��P��9�?�1$0��?}��O���?833333�?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?��X���?l۶m۶�?�r/js�?]t�E]�?���Q� @=��a��?}T$;f)�?�|��O�?�UO���?��(\��@EtA%�?/���}�?�f�M��?��¯�D�?���Q�@%�����?*��RJ)@f|��O�?D0��fa�?�G�z�?�m�=���?WUUUU��?���a�?v{�e��?���Q��?��A!K��?r�q��?�=�� �?�١�?�G�z
@����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?��״��?Ѻ���@��O��?����T�?���(\��?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?_^MiK��?�q�q�?P����?@�wܛ+�?\���(\�?)�x�?UUUUUU�?JB��EX�?�-�t�b�?q=
ףp@�t�!O�?��+��+�?��\�2�?�2����?`���(\�?����?CBq�n�?�M���?ABЋf��?hfffff@=B�k��?g�K1_h�?;9�=-�?$�D"��?q=
ףp�?���|�?      �?��`��?iiiiii�?{�G�z@����Z�?+�O��d�?���s�?���rD��?������@�|��	�?b�־a�?pA�D�?���rȔ�?H�z�G@����Z�?r��Z�@� ��r�?g��|�Q�?033333�a�B��?�������?' Z�u�?�����?���Q�@P�����?UUUUUU�?�k�1���?O�n�	�?��Q�@Za�T�
�?�1���N�?D��car�?�MҷV��?H�z�G@:N�1��?G�:y�?Y<�&!�?F����?��(\���?�o�����?��%�̀�?�\"�0�?P[AG:��?�(\����?J^��&�?���d�?���w�?�\;0��?������@����?      �?ŵ�a��? )O��?      @�6�)��?7�S\2�?�^�r��?�kD�
��?�G�z�@y��RE�?n,�Ra�?�$\Z�?��S�p�?�������? �	�'��?pN�F��?�^mSz��?�]�P�?�(\����n#�{�?%z�$z��?0�1��k�?��M�<��?      @@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?\��Z�?�$I�$I�?��ԉ#\�?����>4�?]���(\@\�f��p�?� ���?�Z���?�Ytl�?�G�z��?������?������?�X^o�?��<t/�?H�z�G�?4s���?�����?/z�V�4�?~"����?H�z�G�?���[�?����NB�?b%c�r�?����]�?hfffff@�J�LT)�?�������?5�Z(��?XV��?��Q�@�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?h�����?��1����?�IF��?�_{�e��?��G�zĿϙΔ�?a#@i��?M��d�?��,��?      �?evoƃ��?�q�u�?�)���R�?t������?0\���(�?L�Q���?����S��? 0 ��?4և����?433333�?�l���!�?�9�s��?�1�[x}�?�[��"e�?*\���(
@_i�"�?VUUUU��?��i��?)\���(�?�������?t��!���?,�X��?^*��U��?�:�>c�?��Q��@�`�5^��?-iKڒ��?t��}��?Ă�� ��?�(\���
@W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=꿾��S��?��c�0��?k��{<j�?9
�
0�?<
ףp=�?�8s��?�Ox!A��?�Sq#���?/�Ij���?�G�z�@޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?����q��?      �?M��7���?      �?�G�z @KY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(�X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?�
⛏A�?��P���?4 ��<�?(
P�;�?������@��t�j�?��qg	��?d���1�?(�)��;�?�������?�T����?Z7�"�u@m�����?����T�?�������?���1�?��fy��?���N�R�?Wŵ.���?���(\�@���n��?�n0E>�?T3	Z�e�?xH����?R���Q
@�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�W���?{�n��?	sG�h��?в�9��?��(\���?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?[��`��?ك2�*j�?� �;��?�������?�(\����?P,��v�?�������?4:�$�x�?�%����?�G�z�?��*�?9�&oe�?ߘ�[]�?��Я[[�?��(\��@y�-[Y�?�8�?'�8����?%���E�?�G�z�@������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z������?�N̓���?�[����?*) �'�?\���(\	@�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?G���;�?�x+�R�?gj��?�r4.G��?��Q�@J��YL�?VUUUUU�?!��a���?�7�7�7�?      @�ao�2 �?�Λ�~b�?����?H݊ÿ�?���(\�ҿT,���?T:�g *�?"�[��t�?7.Hj��?�������??d~-��?�u�����?����2�?� ?7��?      �?E�X9�x�?-��,�?)=��'�?��0���?�Q����?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?{��*W��?     @�E!��p�?�$I�$��?�G�z��?�ݭ����?yþ�\�?�CM`��?�w��K�?�p=
��?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?�r�>J�?�|���?n1DE-[�?|�,����?�z�G�@�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@@>`]p�?;�;��?�����?���O��?������
@�O�<�?������@uq_�E�?��$2��?H�z�G�?����em�?׊��+��?Y�����?"$�A���?�(\���@�83���?�{Nm{�?�F�� �?�������?P���Q�?��0��?R�}�=�?ӗYl�n�?.�袋.�?�Q���@}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@3�J���?�F�tj�?^���i��?�
� ��?�Q����?�D�;$�?���&�?�p߃���?��N�M�?�G�z@��K_`�?      �?��]�q�?�eP*L��?R���Q@�'���?�*H^�?�����?Oozӛ��?,\���(�?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?�S�����?���NV��?��=��?^���?��Q�@P5��3*�?Y�eY�e�?/�G�a�?�M6�d��?H�z�G@
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�������?�$I�$I@��;���?R���Q�?�z�G��?N"����?FFFFFF�?�-5��?����o�?��(\��@뀂���?��Bt�?�(�=l�?��ұ�?أp=
�	@Po�S3�?!1ogH��?�8Sn�Z�?8Q�H��?�Q���@!��m#�?r�q��?�_پ%T�?"Y�B�?{�G�z@M؜�ƹ�?x�5?,�?a�}�I<�?��Z%��?��Q��@T-����?UUUUUU�?L�5���?�������?ffffff @փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?�o��5�?O�o���?�7��ֲ�?J"���?�(\���@����0��?�x��ܷ�?Y1"�	l�?l#֥���?��Q��	@�n���?H���x�?6?�x�o�?�#�	<�?R���Q@�'=��?��fě�?��Xf[�?���¯��?�G�z @6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?Q�����?I�$I�$�?���Y�?z��!y�?333333�?�@����?�����?���Q{�?(������?�p=
ף@5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?��� ��?:��8���?��'c��?�-Wr�?333333@�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?��S3;��?ĸ_�T>�?��a8%��?�,�י��?q=
ףp@�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�_����?      @����,��?[�o�W��?���Q��?8P��A��?�\;0��?<b���e�?y{�X�?      �?~�W�f��?y@�z��?�{b�?�W�^�z�?�z�G�@I��q��?�'iq��?�&��?#�����?�Q����?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?0	�`���?o�vu�?N�� V�?��X���?��Q���?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?���RG��?"�u�)��?��s��?��o����?�z�G��?Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿ�h�(���?����?�3��=�?g�=���?�������?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?��n9�
�?�Zg_D��?_j�P�?r1Bm��?H�z�G@lq�����?ѭ8��7�?�V8Y+��?��07�Z�?������ܿB���?������?��yk�f�?|��¬F�?�Q���@��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?_�;I*��?k��FX�?e�5���?J����?R���Q@�d����?���-���?_l�9��?L��N���?P���Q�?�{����?�Pd����?�{c����?�������?���(\��?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�?�}�!���?��Sڃ�?xE.�;	�?��}A�?��Q�@�]�L�b�?2&�l�?      �?]|�c���?�z�G�@�va�q�?iiiiii@�;��`�?      �?433333�?P��-��?�NV�#�?8��m���?�;�#�?333333@�G,���?�	����?���R{�?��?�c��?���Q��?G�u���?�t��6�?ZM��W�?�ɵ��?gfffff@{^Q�h�?       @��Tf,�?�7�7�?�G�z @�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?Sª����?      �?�	*�/�?W�<�?R���Q@5~�lk��?u32"��?8����j�?�����?�z�G��?��Sr��?U����?<����?w�{��?<
ףp=�?��aJ��?��˝��?�D�y�?�$���?���(\� @u�-BK�?��T��K�?��x���?>���~��?���Q��?e�Y���?(������?�[����?������?��Q���?�q� .�?��"E��?�V���2�?�^�^�?�G�z�?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?��]���?[�[�@�{�q�?.q����?���Q��?}9�ot��?d����.�?֐��<�?OP�?�z�G��?%���y��?a8B��?�!!?�Z�?���q6�?<
ףp=�?��]��S�?�z�����?����?1�0��?(\���(�?��E4�?Dio����?J_��_�?�����?      @� �����?{ӛ����?��*��I�?"�nd=6�?������@ ��2�?S�n0�?���&�_�?I%�e��?�������?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?Ũ���?WUUUUU�?%�[P�~�?�������?�(\���@�m�02��?;r����?���	���?����<�?��(\���?"ۼ7@��?�q�q�?=ȋ��?H�z�G�?{�G�z�?�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?�{㘺�?zR}%��?!�yV^�?��ծm4�?�(\���@����t�?���j?�?��y��X�?sƎ�e�?������@E� �?      �?��ԉj��?��|�nS�?333333	@��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?|A� *��?�袋.�@��k{�?W�+���?H�z�G�?��r���?\��[���?�4�.��?2}~k���?��Q���?��1���?wF]�K��?={��?������?�Q����?���X �?�\�\�?6#�|a�?>6:8���?P���Q�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?��;��?*b�����?�0����?�8+?!��?���Q�
@� �����?r�q��?܌��! �?���[���?��Q��ۿ,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp��j�с�?�dn}�?�xJ�Rn�?��寖�?�z�G�@X���A�?������ @<�z^��?C���,�?�������?(tҶ��?�/�I��?lv��7��?��cy���?      @��n �\�?�q�q�?!��s �?5/�D�)�?�p=
ף@��{G�?����S�?Y�_��?�����B�?֣p=
��?��mW(��?333333�?"�*|��?���?333333@��[�à�?��b����?��y�xi�?�cp>��?�z�G��?��wW�?�.�E��?K^�3v�?�������?�G�z@�!ފ�?c����?��J%%�?��(\���?�G�z�?]��{��?�����?Iy���?E�,V!�?�Q���@h��Ƅ��?UUUUUU�?���t�?     ��?q=
ףp@�,��o*�?���tT�?Eg���?�@i�
�?��������S;>���?�Y���?�gS���?U�j�o�?أp=
��?P�H �?:��8���?Ta�z`�?�'�����?�G�z�@�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?əPB�?��.���?gL0�h�?l��(�?ףp=
�?V�gb�?��W�l��?U�����?_�HI��?�������?��B~���?ƶ#e��?-��k4�??&ǒ::�?{�G�z@�L���z�?X�O���?��F�{�?!���c��?�(\����?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��<���?      �?��(�r�?��a	G��?���(\�@��m��?����?&z`�5�?2u�=�S�?      �?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?"&�H
�?�?�4��yO�?��)��?
ףp=
�?[�_�?r���&T�?Vl;!t��?�O��O��?�Q���?u��=M	�?�ڧΪu�?f>����?: 2ܫ`�?�p=
ף�?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?v��� �?o}$�o<�?��(ET��?�{i�"8�?���Q�
@~�aE�?"�z\��?�R����?I��/�?.\���(�?ӏK�K�?��{���?���S��?{���g�?P���Q�?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�`���`��?���-��?����w�?��-�jL�?��(\��ſwJ��L��?S��?�p���?�������?
ףp=
@�X��S��?      �?Ѹ�U�?1�0��?���Q��������?�Qf�,�?z�<���?�%���x�?Z���(\@r>bܘ�?��MmjS�?e�����?|1����?���(\��?��B\&�?�n0E>��?���L�?2 K��?�(\����?[̽e��?�)`>�]�?i���/��?o��[�?������?q�ک��?      @���<X�?��=���?333333�?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?�uf�K��?EDDDDD�?ޮ@l�Q�?�������?      @n,���$�?����b)�?A�쎑��?@�1���?
ףp=
@����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?�_�^�/�?      �?K��>�?0�9�a�?������@P@��}�?��k���?      �?�J���?�������?���+*�?�-шs��?���ҋ�?�#o��?q=
ףp@���fR�?:�:��?�Pk����?ק�����?��Q�	@�+����?�#�;��?��oa��?��8���?�Q���ѿΛ��e.�?�{a���?�D1[�U�?Z��Y���?�z�G�@�miV���?�U�;���?P�l�V��?A�Iݗ�?�z�G�@_������?���h��?�����?\t�E]�?�������?Y/�7�/�?�>�J�?��	���?t�����?���Q�@���]�?��g����?1sJJ��?��f$/��?���Q�@\������?���J���?�9�߀�?n/�d��?��Q��@F��W~�?��f=Q��?�����?DDDDDD�?P���Q�?�]A6�?��0�:�?A�B)���?7��O	�?�G�z@A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?*����?{���\�?�N�ҝ�?�����?�Q���	@XD"���?R��+Q�?$ ����?�#F���?P���Q@��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?����g��?�]����?P�øW�?v�=H]��?��Q���?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?auȒ���?�v%jW�@��s5��?`����?�Q����?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?�74J�_�?*6\u��?�$8����?�/t���?      @����?���a���?Û�P�?�`8wC�?P���Q�?�p�|���?���)��?^�3���?h�J� :�?�Q����?l,����?gH���?���2G�?v�A����?�z�G��?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?����?��R�y�?�����?�s@ڦ�?�p=
ף�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?������?�~H���?U��oW�?��S�r
�?
ףp=
�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?������?�5��P^�?lN�b�Y�?���v�?�G�z�@D���Oz�?PuPu�?      �?٫��J�?���Q��?������?�N��N��?��U>R
�?	f���?�G�z@�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?W����?��8��8�?      �?Au���?�������?lv��?*.�u��?m�����?O�<�"�?!��Q��?��i�,�?ףp=
��?���b��?,Fڱ�?��Q�@�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?L�|9��?m���X��?�B�q��?����:.�?833333�?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?�c��)�?c��4�?�.fxx�?�Ŗ����?������@�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿ,"�j�%�?,-----�?'狗�8�?�`�����?133333�?�wF�?��D'�?6������?�_�_�?�������?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ�N"H��?����?Hx`2��?��r:���?������@�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff��
�&af-�??�?��?�q-���?��	�{�?أp=
��?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ�4����?�%����?�J:��?v{�e��?���(\��?Z�yv�<�?��a�
��?��ࣹO�?:&߭��?��Q��@�מ���?�i�i�?Q�XW��?�R�~���?      �?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?��,���?�z�G��?����U��?a���{�?      �?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?��j�G�?u�5�o��?���d��?�~��?�G�z��?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@2�7���?���A�?���i���?_7��T�?R���Q@c&i�?�ÔP��?P>�z��?�uI�ø�?      �?+e��R�?pА����?�_P�
�?���譺�?��(\����܎h�?��/�$�?�p\��?���6�?���(\��?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?��I��?      �?	)�L��?ڟ�!T�?��G�z����#���?�rcˍ-�?���'��?8��{�?@�z�G�?(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?��=O�?M4�DM�?���2��?�ܛ���?
ףp=
@@�X兞�?f���?����15�?�>��?��Q���?erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?O�TE���?�(፦@��x�b�?��RJ)��?�������?f��UJ��?�!XG��?�����?����vW�?8
ףp=�mӞ��?#��~j��?�1?��l�?��i���?�Q����?��zZ �?&jW�v%�?t���?X`��?!��Q��?;�H�r��?W�rCH�?��A�^�?�����?(\���(�?	�F@�?�����?c�I���?l��&�l�?!��Q��?����*�?)#�`��?��@�x�?�gL���?أp=
�@:����?�5��P�?v$����?;�;��?أp=
��?9gήc��?�Z$�R��?������?�/��/��?033333�6%�M���?���s @N�|ҍV�?e�e��?�������?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?��X��?�Kh/��?�f i5�?*g���?���Q��?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�n��?�3_�g��?����B�?`V�4[s�?`fffff����/����?���T4�?h�v�Q�?�����? ףp=
�� '�Q�^�?ᖚ�?C�7�y�?4H�4H��?���(\�@
��Y0�?�G*;�?      �?������?��Q��?/������?�k��%�?���g���?8S����?�G�z���뚖f�?1ܫ`���?��Z(~�?�;�;�?@\���(̿�����?�DxR���?`f�"�?�8yh=�?q=
ףp�?��
�?�"nps�?�`>J�?/������?���(\�ҿ���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?qCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�  I   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM�qPh"�Bp  ?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����?P����'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@M�4i�@'M�4i�@'M�4i�@'M�4i�@'M�4i�@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�C���X��?qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�CeC���9�?q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�C����6W��qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�C���X��qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM�qvh"�Bp  ?P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����??P����?'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��'M�4i��M�4i��'M�4i��'M�4i��'M�4i��'M�4i��qwtqxbX   _sklearn_versionqyX   0.21.3qzub.