�csklearn.svm._classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX
   break_tiesq�X   kernelqX   rbfqX   degreeqKX   gammaq	G?PbM���X   coef0q
G        X   tolqG?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq�X   max_iterqJ����X   random_stateqKXX   _sparseq�X   n_features_in_qKX   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
q X   f8q!K K�q"Rq#(KX   <q$NNNJ����J����K tq%b�C      �?      �?q&tq'bX   classes_q(hhK �q)h�q*Rq+(KK�q,h X   i8q-K K�q.Rq/(Kh$NNNJ����J����K tq0b�C               q1tq2bX   _gammaq3G?PbM���X   support_q4hhK �q5h�q6Rq7(KMM�q8h X   i4q9K K�q:Rq;(Kh$NNNJ����J����K tq<b�B4	                                                   !   #   &   '   +   .   /   1   4   5   7   8   :   >   @   A   B   C   F   G   I   J   L   M   Q   S   T   U   W   Z   [   ^   _   `   c   d   e   h   i   j   k   l   p   u   v   z   |   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                !  "  $  &  (  *  +  ,  1  3  5  7  9  <  =  >  A  C  D  F  G  H  K  O  R  T  U  V  W  X  Y  [  `  b  c  d  g  h  k  l  m  p  q  s  t  u  w  y  z  {  |  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                                   !  "  %  )  +  .  0  3  4  5  8  9  >  ?  @  B  C  D  E  H  J  N  Q  R  U  V  W  Y         6   P   Y   a   g   n   w   �   �   �   �   �   �   �   �     -  ;  I  S  Z  e  }  �  �  �  �        #  (  ,  /  2  7  F  [  \  ]  ^  k  l  m  n  q  r  s  t  u  v  w  z  {  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �       	                       !  "  #  $  %  &  '  (  +  ,  -  .  /  0  1  2  3  4  5  6  7  8  9  :  ;  <  =  >  ?  @  A  B  C  L  M  N  O  P  Q  R  S  T  [  \  ]  ^  _  `  a  b  c  d  e  f  g  h  n  p  u  z  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �      q=tq>bX   support_vectors_q?hhK �q@h�qARqB(KMMK�qCh#�Bpn  �h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?!}u�O5�?��=Qr�?7r#7r#�?y�sJiM�? ��c��?433333�?�Qa���?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��?aC�����?     �?J�.����?"1ogH��?��(\���?|UKP�_�?
��Y0�?�G*;�?      �?������?��Q��?�-�����?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?鄣Z��?��״��?Ѻ���@��O��?����T�?���(\��?���7 g�?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�z����?�!ފ�?c����?��J%%�?��(\���?�G�z�?�~���?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?f��UJ��?�!XG��?�����?����vW�?8
ףp=��,���?p;̞��?      @�њ�%g�?'u_[�?�������?y�l��?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?עWG�?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?r6]����?�������?�	��6f�?���3$��?H�z�G@��S��?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?���. �?i�`���@jڪ���?��}ylE�?�(\����?ڔ��ɣ�?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?�a+� �?O9:����?�f^w�O�?y��x���?أp=
��?R��i��?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��K�?�&�j��?7��P^C�?F�����?q=
ףp�?��G�z�?:�5+�?����g��?�]����?P�øW�?v�=H]��?��Q���?-s��ǟ�?�X�y"��?%'¸Lr�?c�/�]�?,mG8��?�G�z��?�^���?Un����?�������?#�R���?]�����?�Q������j;����?��h�D��?��P��9�?�1$0��?}��O���?833333�?&~��.w�?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?��L�F��?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?��2MK�?�`�`�?{���K�?�.�|��?��(\���?�٤�I��?�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�i\|��?Ե7�rL�?�l��l��?���'��?��E���?��G�z��Ψ}Ri�?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?�9vZC��?X7�"�u�?A ��X�?ƃ'��?�G�z�@��n���?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?\	# ���?�߈��?Ľ9�X�?и[���?\���(\�?b�����?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?ű�r��?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�!�/�?P@��}�?��k���?      �?�J���?�������?"t�I�+�?����?��R�y�?�����?�s@ڦ�?�p=
ף�?7���M�?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��?9gήc��?�Z$�R��?������?�/��/��?033333�EF��DG�?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?��[y��?�Ў�e��?��^*)�?z^{�?�(\����?�9)�?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?��O�V�?�m�02��?;r����?���	���?����<�?��(\���?�ca�M��?���?�m۶m�@��X)�O�?�\.�?)\���(�?^�)�Ҝ�?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,�����?�h��g��?O ���E�?��mQx��?��vY��?���(\��?`���+��?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?[�>���?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?It���?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?u��׿�?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@c-�Gb�?�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=��_��#�?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?L�|9��?m���X��?�B�q��?����:.�?833333�?����?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?�M�2�?z&�����?�H(m���?��K�y�?���cY��?��Q���?��ʦ���?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?R8�u�?S{���?��,�1�?:�oO�$�? �G�z��S�hz���?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?��.����?��Sr��?U����?<����?w�{��?<
ףp=�?�c��o�?���~�?9"�P9�?<O�����?!������?���(\��?�c��D��?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?�'=��?��fě�?��Xf[�?���¯��?�G�z @���#��?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?{��*W��?     @�E!��p�?�$I�$��?�G�z��?�_�����?c�2��8�?l�l��?�����?T��S���?�p=
ף�? ���P��?���g
�?&���^B@���X^�?��FS���?G�z�G�?;��q�?�D̥�
�?�Zk����?��iz�?���\��?��Q���?��е:�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?�՜�pH�?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?U@�'��?�x+�R�??dM2_�?�(S�\��?�(\����B��e��?X���A�?������ @<�z^��?C���,�?�������?\��陌�?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff��7�z�<}�?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?      �?���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?�'LZ��?���e��?I��/�?i�(�U�?�VC��?T���Q�?�74��q�?"
c���?�[�[�?��
y3�?q�M����?���Q��?�����?փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?����y�?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?���#�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�Ǔ���?q�ک��?      @���<X�?��=���?333333�?b�-ч�?��m��?����?&z`�5�?2u�=�S�?      �?��]�E�?ƪ+�K�?~r!�f�?�`(vo��?l��';�?�������? !�!���?�s[W��?�7�P�?Eo�h=�?�r(w��?���(\��?�TS�Yd�?�Ĭ~��?��Q���?>s=��^�?�����?�(\����?�a��~�?,"�j�%�?,-----�?'狗�8�?�`�����?133333�?̕x�F�??d~-��?�u�����?����2�?� ?7��?      �?��Ld��?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?*��Al��?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?i�+s�?333333�?`�>��R�?��.���?q=
ףp@=�f{?��?�מ���?�i�i�?Q�XW��?�R�~���?      �?t��3��?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?ѳ!s��?g�\���?�����?��񍔎�?����.��?�G�z�?'�����?�2�j���?     �?u�;�F�?�$I�$I�?�z�G��?Ud���|�??V�)��?_�_��?      �?��B�
�?�G�z�?�Z�K9��?�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿�_�Be�?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?���+��?��p����?      �?��e�N�?�������?R���Q@>����?(� .b��?�k�S��?��F����?���w���? �G�z�?�&ɢ�X�?�O�<�?������@uq_�E�?��$2��?H�z�G�?aq8���?��aJ��?��˝��?�D�y�?�$���?���(\� @��p��A�?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?`���`��?���-��?����w�?��-�jL�?��(\��ſ�E]�?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?�h�(���?����?�3��=�?g�=���?�������?���w ��?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?�L���z�?X�O���?��F�{�?!���c��?�(\����?�g����?Шx�?jF���?������?�.�?��?�z�G��?��2}��?F��W~�?��f=Q��?�����?DDDDDD�?P���Q�?.����"�?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ʞ2����?��	��?�jL�*�?�\�K	)�?U��t>�?�������?�ϗg�?�ӄ���?R���Q@���K���?����*��?�(\����?I^J��?�
�����?���!y�?��S��?�����?������ܿ����c��?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?6K�b0�?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?9�IA�?����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?]T�%,u�?%n����?      �?7��S�?��/���?�p=
ף@�N�w��?5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?����?�T����?Z7�"�u@m�����?����T�?�������?���ux�?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?_������?���h��?�����?\t�E]�?�������?LkCJ[�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?���-��?�������?�p߃���?y����?hfffff�?fd-c��?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?���/�?톘��=�?+P�W
��?���gk�?�������?Z���(\�?�Q�rX��?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?9�m�.�?�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?#��3�U�?^���O�?o��o��@�H<�'�?�X�%��?�������?�8�T/�?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?�v���?U�����?����?�M����?�(\����?2�g2��?[��`��?ك2�*j�?� �;��?�������?�(\����?,evp��?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?�-{X�?��{�A�?,˲,˲@�Z�rf�?c��0u��?���Q��?��v��?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?J""}��?����;�?jZ��m�?�0�9��?��Q���?Zf����?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�Y��.�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�?u�-BK�?��T��K�?��x���?>���~��?���Q��?f[t��?U[G[��?;�;��?�	v�o�?�a�a�?������@U��A��?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?O�TE���?�(፦@��x�b�?��RJ)��?�������??3�/D�?�_����?��.��@�ʌ����?�v���?��Q���?> �xka�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?��<���?      �?��(�r�?��a	G��?���(\�@n.>��	�?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?�Gq���?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?��zZ �?&jW�v%�?t���?X`��?!��Q��?���f �?�п�cX�?���؜��?��{�z��?�F��?_fffff�?�F�9���?fo/���?/����?'N`�4��?��3���?�������:T�+���?����?      �?ŵ�a��? )O��?      @�����?
��\���?��\AL��?)us�?      �?433333�?@�����?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?+e��R�?pА����?�_P�
�?���譺�?��(\�����f��?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?��9k��?5�T3�?233333@牫;X]�?�������?333333�?��W7�?�i����?T����|�?�;x�]z�?,d!Y��?P���Q�?���}�I�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?���1�^�?C�oB��?      �??��(b-�?b�1`�?433333@��
�f�?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�? ����?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?|A� *��?�袋.�@��k{�?W�+���?H�z�G�?��J.�?�C����?�������?A�ra���?�@۽U��?���Q��?�/�����?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?�~�A
�?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?l�ģC�?/9(��?.�袋.
@�*����?�������?�������?�/%Ŷ��?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp�\��E�%�?�5���?@7���$�?h/�����?�������?�y;Cb�?s��&�?(W�7�?���xW�?B�HV��?��(\���?�LGuk�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?��F�#�?�Q���?������
@>���fi�?_*�-5�?�z�G��?� +\�?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?6%�M���?���s @N�|ҍV�?e�e��?�������?�� ��?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?m.���?Q^Cy�@��=,��?_�ڕ�]�?\���(\�?���^y�?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�? ��2�?S�n0�?���&�_�?I%�e��?�������?����5�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�9��-c�?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�<�^�?"K�_y�?���,d�?���<�?jhɬ�?�Q���?D�&Dq�?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���?P,��v�?�������?4:�$�x�?�%����?�G�z�?Qj����?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?:r����?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�m�����?�X$����?L�:,��?&����?G�N��?\���(�?�'�	�?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?'���/��?��
�	�?:[���:�?�!!?�Z�?�0݂k��?�p=
ף�?̓�lXD�? �5�0��?�����?B �Gey�?r�q��?��Q���?���I���?ϙΔ�?a#@i��?M��d�?��,��?      �?;���?I��q��?�'iq��?�&��?#�����?�Q����?�E��Q�?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?K]E!�6�?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?=������?��f���?O���7h�?���t��?���(\��?՛>����?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�vף]��?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�??4G0�?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?m��C�?      �?2zW�]6�?��L��?���(\�@��y����?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ(�~��?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�??[�w(�?�>����?      �?0`z��Q�?'u_�?�p=
ף�?W�n��~�?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?�a��P�?����/��?~�~��?LgR�L��?|huq���?�p=
ף�?�8G��s�?�N"H��?����?Hx`2��?��r:���?������@�P	�_�?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?�{����?�Pd����?�{c����?�������?���(\��?�ֺ��	�?��9���?�e���?��G��\�?�����\�?���(\��?:����?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?*����Z�?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�b=��
�?<�b���?����?�Pp���?Ŕ��%�?�p=
ף�?�����?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?vP�I��?E8S8B�?������?�5��P^�?����������(�?��I��?      �?	)�L��?ڟ�!T�?��G�z����8I;�?�G,���?�	����?���R{�?��?�c��?���Q��?;⟯�:�?}9�ot��?d����.�?֐��<�?OP�?�z�G��?�dn�>�?��B\&�?�n0E>��?���L�?2 K��?�(\����?O(���?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?T�.�n��?�-�׮�?H{����?������?P���Q�?��/>�?�܎h�?��/�$�?�p\��?���6�?���(\��?�=
��y�?:����?�5��P�?v$����?;�;��?أp=
��?�[9�.�?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?���A��?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?Xe�6�?
ףp=
@�3��x�?�D�Z���?(\���(�?2�b���?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�w�x@�?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?P�ϸ=�?�YĘ��?9��8���?�鑢3�?^��3��?�G�z��?�*ml|��?��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�?����j��?auȒ���?�v%jW�@��s5��?`����?�Q����?��LO��?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@yU�٬�?�83���?�{Nm{�?�F�� �?�������?P���Q�?1l(�?e�F-��?�������?���:%�?V���g�?ףp=
�?´�z�)�?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?lv��?*.�u��?m�����?O�<�"�?!��Q��?��P�)�?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?֊�q��?��Z��Z@�K��?#e�����?���Q��?
k#w��?J��:���?=
ףp=@��=!E�?���E�?=
ףp=�?O����?��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?�?w�q �?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�`1+�H�?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?��X��?�Kh/��?�f i5�?*g���?���Q��?{V�|4�?�,B�N�?�
��v��?�߾���?������?P���Q�?z��V��?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?^` 5��?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��A��?�P�6Ԗ�?s>�cp�?�`κ��?���$D�?P���Q�?爈��P�?���\�?�^o�?�?Q�/��?^̧^̧�?�(\����?�XrYǾ�?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?�X��e�?q����?*�3��?3iM��h�?QJ)��R�?=
ףp=�?��U#3��?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?V�gb�?��W�l��?U�����?_�HI��?�������?��h~3�?F}�p �?������?N6����?\����?ffffff�?�T����?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?�S�����?8�P\�?��;^�?M�*g��?\���(\�?�	�;D�?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�<��2��?2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�V����?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?�
>U�?
ŭP�
�?Pf�i���? i]���?�G�z��?�_����?���;��?���˦�?Q
�C�?����1�?�G�z�?��1�2�?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?��j�G�?u�5�o��?���d��?�~��?�G�z��?\�o�nl�?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?���q&��?      �?�ƽ7�?%Ԑ�W��?�z�G��?4�^}9�?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�	ږ@��?�3��j5�?l�O����?�4`Zz�?n�s�p5�?H�z�G�?5�H���?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@��Y���?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?v�����?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�����?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�s����?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?t��Y��?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?M\=���?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�\��f��?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?|? ��@�?�q� .�?��"E��?�V���2�?�^�^�?�G�z�?Hݽr�?gDAl���?<e�U!�?��-��?'u_[�?�Q����?"�R[WD�?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?�_{��\�?�S�����?���NV��?��=��?^���?��Q�@�D�y*��?�������?�m����?G��|���?E4Z����?�z�G��?hE�-\�?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?���p9�? Jx5��?�a�a�?�;x��<�?�������?�Q���@8)���>�?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?���V��?�'���?�*H^�?�����?Oozӛ��?,\���(�?��x~q��?�wF�?��D'�?6������?�_�_�?�������?�Ko��?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?:��]��?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��76�?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?g?�V.�?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?���6���?�w���?zkfkl��?�k(���?      @�q�^��?"�FU��?�71}�?v��3���?�N�Q�S�?�Q����?�5�,[�?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?Ŝ�lK�?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�X�!)b�?X�!c��?���a0��?$��P�?���'a�?�e�<O#�?����v%�?)J���?ڇ��y��?�v	�2�?b��Kw�?~Px�A�?�'���?�/'�(��?:Q�}��?O���2�?M]�=���?�/����?n�����?����u�?@R vr��?��5��)�?;B�^Y
�?�";cs�?ɮ��0��?�}T��"�?S�S��?������?��c����?�A�2���?�X�*��?��ȱ�?�5��\�??V��?�kgea�?�UAg��?����2�?��^���?˶��;�?��EqFu�?�Q{wpA�?�YH�4r�?����c�?9^�N��?��/!�?�t��b��?hm�)��?�ګ��?ky�/���?nM^f>�?i�`���?م�Y�y�?�,|�?6��R��?9�.A���?�'�6�[�?�a�>�E�?~2�㶂�?�x ��w�?.������?�Z�հ�?p �&?�?���o;T�?\Txk��?���m�?���+̀�?c"X4` �?�jM I�?T�ΗJ��?շ�R&y�?t�۽���?8�;���?ɶᰪ�?��WY_�?y�Ke1�?$崪+u�?5$f�Г�?�	:�S��?�{���i�?�V7�FC�?�%2fm�?lY��y�?jؙ�T�?���t�#�?��]���?]}�BC�?) Ld[��?q<�
�u�?��iz��?:c��3�?A�-��Y�?vcutT�?�ٌ4l�?aN��?,e-v�?�~����?9�V�q��?e^��M��?�y3ʆ��?�*��b�?���:-�?���~�f�?��uv�?�e.!ݸ�?�"*ͫj�?�P�>g�?�PH���?�T}.��?H�'}��?px�� �?b�2w��?4C_N��?/��D�?�U�b�a�?��E���?3�"���?��V����?���W��?����?�t�SK�?�L�i��? �т��?����~8�?7:�*�o�?ё�:%%�?����"�?�>���?Wr�ݭ�?BҨc��?��l��?g�����?`�׌j��?�;�]�*�?~XЧ��?I���r#�?z���Es�?��?�#�?�NCߵn�?��c�e��?�����?:�.C�?ʁT7��?#�-Ɂ��?����c�?׳kA�?֌{7� �?�}s�J<�?.��#���?c�_F��?�������?�a�<j"�?H���X�?�'fپ��?J�#�?˴;�ah�?���6��?�=�c�	�?�"8��?�_ЕI\�?2J���?�s�J�y�?�VХO�?Ճ�$��?<�ĳ�?O����?`�~���?|Ga�L�?j��p�r�?J���mK�?5$��2"�?����U��?�aT�? �tC�5�?���%��?�����?"�N)x�?�c+��.�?�5xn��?">ZNf�?l��Ol�@�p��X-�?��(͆�?<�Ey�%�?����;�?�X3 �o�?y
�a5@��D��
�?~��\�?.��a��?�++��?�33�w�?0���@a=���r�?eE[���?L���qu�?�!�G.�?���޶�?�s8�
�@���D��?(P�K�2�?�v���?h�V��/�?�˲7)�?p�.�@Nl��d�?{���'�?��E��?��q4�?n��Q)E�?�TI��@R���?d} v�%�?rӈ��?���M�?g������?Ha��� @��@Ɍ\�?��X�ey�?Yx��m��?�i�AN�?1���>�?�jS?�?�g@�X�?9�I�`��?]�o��?EO�l�2�?�^���?�U�\q�?y.�h��?vr} W�?2��.��?�h�`�%�?�-c��7�?��e��@��X����?cT����?a���'�?�'��9�?��Y?���?c�F���?���^2��?'c�=��?���]��?jеXj��?/0i����?�R���@�`��%�?�g��O��?�����?��o0�?\����v�?bڐlT[�?�f�ܙ��?��!��?*��#}T�?Ұ��@��?H�I����?}���,^@ͧM�}�?��w���?T�z�k�?i%;5���?"����r�?k��`b�?���~�?���R�l�?�H3*��?��{\(�?ߔ�}>�?nx����?fF�W��?�Eb���?�<�R���?�~���?o1FJ�=�?-2|�0�?睃vɉ�?	��9��?&�Ϻ���?U��?G��ΠI�?�"��T�?�B�+��?nq���?aF����?�$3�N��?�)�$:�?��F���?q�mMm�?c�1��y�?c�Er�?`��#��?� =4
�?_�b��?����?�mr1�;�?3d���?H9�����?Br�)�?׫�`N�?\ ?��?��rݗ�?U�;�(�?�Gr1�?W��sp�?�!��@�?��|)�?[:����?�w��4R @�wRl��?$�k��)�?"����C�? 2P&p��?�B_��?\9: �5 @�h�y��?�bjk��?�)x�;�?�)#��?�o(�^�?����#��?<n�r��?�'n�?�?W�aVj|�?v�w,�V�?d��ww�?h5�""+�?�o)�w��?�U�AN�?<�OIN�@N�֌d\�?ÁC��1�?HiM��?�^��/�?[���+�?�)η@��dR�r�?H3� m�?�ۜj�Z�?<fV̓*�?a�(p���?�³�~@�&ty���?�\L,��?8�s�lb�?��֑P�?�r�s!��?�c��xR@W�w�?��(a���?��t��o�?9�"U�?
n��m�?��<Eb @ �`w��?8��{�#�?H�+��?��6�?�t鮅N�?�8-!u@(q���H�?L����O�?���G���?���}��?�\�����?�M�6@���m��?V~��?�H����?��R��8�?�51^�?��HW@��MhШ�?�h��d�?q$�"9�?Ynh�(�?���I���?1Q���@P/8��?�͕f��?m�����?�Y�Vw�?�2�y��?�	�s��?���<��?<��#��?(�mw���?�5R�v�?�\'���?��뿊��?杠���?Q���R�?�f��s��?�E�$h��?k�D�7�?��{�̡�?��b�D��?�nRjD�?��5È4�?�7Fw���?f���3�? m���?ݞ��y�?.�lD�?�^�.�]�?%�xfޚ�?���,�
�?����y�?�R ���?Q]`�5�?5}�0���?�����?�Z)���?ƕ��Q�?��5��?x
��>J�?$�SNͩ�?��F���?A��ؽ�?�otƂ�?N�]�?i������? ˘����?I(kc^�?���- h�?l,�어�?�.N�#�?�][[Dw�?�F�V��?����O�?	m�q8G�?�E�u��?3m�ZA�?���o��?#U�34<�?��X�/3�?H!�N���?$���b��?�����?�L-2��?�5|V�B�?Kbg>[B�?��"��=�?N'Z�{/�?�ډ���?L��Ӑ��?2�Ż5�?��~�b�?p���9��?�Sݐg� @#��Q�3�?Z���y��?l<����?u��Y�P�?	�"�p�?*�����?�5v!G��?�o����?����O�?	:�x�b�?�͛�|�?L��=d1@(w7�b��?�ح{��?ɔu��8�?Hc�?�S�uw�?z��K�;@��X���?m�(��?uG�
)��?����BI�?|O�U�?tVX-���?Otr_]O�?�U�^�!�?�n���j�??mFұ�?l�#.���?ɷw,+�?Ke���+�?�]�� �?�f=�o��?o`����?F�Q��?F*_OA�?�$�=�R�?y�{g��?�^��/�?s��m���?:z.�q�?�c&Qs�?T�ʼ@��?�V��>�?�NRAN��?����?on���?�
/�"�?lΗ�t�?�C�����?˜�V��?z�K'���?���c��?bq9���?�oaA�-�?�#����?О���?;W4����? ,x��? ��Ā��?F{�PS��?'������?���?���?��oS���?H����?�����?E�Y�9�?�9�W��?"�-cZR�?|���@j�?��·X�?*���?h����?�������?n�>��U�?��VY�?��i���?L�V�?�)/�?��ÎV��?~#��5��?���W�?G�)�y��?�M���?�V�Y��?��}Ǖ��?y���b��?�?��U�?����?L�{�K��?�;$.V��?!t��
�?���.Z{�?=?t_���?o�{���?���p�?n/� �J�?=x�?N��5�?0]��R��?����s;�?
���F��?,�=�O��?�*�U��?)]�Wj��?�0r\��?f�b���?9�ur�V�?(���L��?E̲#�?���f���?�W:%���?����g�?Y؆3��?��13~�?2�oǜM�?!!��H@��k�?�x�Pf��?���W�?���of�?�����?�?���`c@��˻n�?�J� *�?~��o��?\�����?��2�#.�?��v�< @�)�I��?�"
5���?�O���?B=���$�?��%�?�e1���?E����?�a#�X�?�H����?
ƒdۮ�?�5����?j�"R @pU<��?�<����?�1�q9>�?�q����?e�ʀ�Q�?�5��v�@vU˯�?��S:h�?0N|��?
K���?���  �?w��@���?W�q�Ή�?ZxR��v�?��mHnE�?���~�?��~���?�z.W�y�?}�:��r�?8�����?��Pb��?8&���?RՊR%�?$Ŗvt��?> 
=��?M�k|��?��hZĭ�?����^�?��f�a�?��t���?!��>��?w=�t���?&p�H�?���t���?��+���?.:wl/�?
S�R��?�K�FɅ�?�=���R�?^]H��8�?���*1�?�7�x��?X������? ���N�?;����?�dA�nU�?��e��?�(��8��?y2cd�?����?�����?���yk�?&�u��%�?6��Vt�?�G*'�?��Is�?db C���?ql1k�?ad���-�?za9�i��?����2�?�J���]�?�9�AB�?d�_�q�?�B.��)�?[��4�-�?a�r�,�?�S���h�?VK�5\�?Bg3��n�?�yDy(�?�yf��?4�-�?�=6�P�?麽����?�U�DG�?.W��+��?�z@�"AB�e�?<��x^�?R���%�?'6�S�?�c'����?�|E��@ R�e>h�?���M�?x�rl���?��bl��?X���{��?��D5sp@&��4Kc�?��X,�l�?��sWT�?A�$)��?����8�?7�F�D��?U�p�l0�?<�sP�?'�bҩ�?��^�T��?���Q��?V{�d��?e�Џ��?�7"i���?�ޮ���@�p�����?Z�����?B�̲��?`�M~T��?ʨ��S�?���C��?���X6R�?��bY	��?�I��z��?� ���?&��暲�?�� |'��?p�����?�L���?�cB4W�?�&O+/�? k~���?�.��@A��qk}�?����ڞ�?nP�?�cP4�?¶�N��?ʱ�$e}�?[cq���?��ۯ��?�g��mz�?Wa�l��?i'@
��?��[8�5 @����I�?��%>���?�w�'�?�������?�01��?`���r��?���;�?���%��?�8����?Of�u��?���'B�?o�F�?�}�1�3�?��_;���?����vO�?���.��?�T
���?W��x�?s<$�?��,���?T���v��?,��,���?������?Ð�C��?��3�?FX���?��+�D�?B�2�H�?�L1چ��?��P��?�k L�?�P?��?t�Ŕf��?$����?�U01���?���=/��?�j,� �?L�?|��?8{���6�?�w�`��?�Fe\O��?����?X�?E����Q�?LNf)�?����в�?<J�(�?r����?ʸ.~+��?��O���?�}�z)�?��a�*J�?C��vܼ�?�08\���?H:�r�?ytʥ�w�?�@\_�-�?�����m�?FZU��?�(q��=�?�mid��?���7�?hs��
�?��v'��?�t����?>Lf����?�/Ȋ�~�?��H�?����'�?�f���?���h��?ޮ.}A �?� ��a�?P�@�t�?>����?W���[�?_bt�\��?SHZ`��?ڂ�U@�C�P��?
����?H���?��s���?�UL�	��?�5ohx4@O�ѿ��?.Ls׾�?��b���?��ߐa��?!v�l��?�Ok<@2�����?��h�W�?�Q�'�?P7c���?�T�ݱ�?��c�m�@��V�"�?Wy�r��?��TA��?
Rg���?JO����?^�Jp1@0��k��?K�`�� �?@��	rr�?���!�?���c��?6���;@�GC"��?e�?:���?��/\��?s"�#{��?Φ�$O��?zvJ��?6�z�[�?q_�,��?h%��?�xc�P��?iC�}��?��A��?yi�,if�?����?H��4%�?3��j}�?g���F�?�D�s���?~dx,N�?Y�2�3�?5��AZ�?�*�w��?�6n��i�?�#'����?><�u*��?,!�5���?0%`/��?���H1Z�?������?�朖r�@���۴��?Yɴr)��?}�3*g�?�Q���<�?�l�oF��?�Pt8��@d��9?�?��?���?r�,���?���V��?��P*��?�Y���@�hJO`�?0r]����?�A��[�?	:����?�H��0�?1$�n�@B?�	��??�Ov��?�g�����?����{��?
��o��?z*"�"�@Fa��@��?��U���?q�3�_��?x:��ϸ�?e!�͡p�?�e]l -�?���x��?O��f��?U�f�7��?�U`���?��T���?�?,�+�?G��$��?�c�t�)�?ʙ�����?,��˥�?�5����?��opQ�?8����K�?Rt��"�?���?�	���?�U�R�?L��"���?b�&�?C���R"�?�9PZ��?�0#���?�&ƘQT�?�������?uzl��?&��i,�?
�����?�C�	���?ۤ�0�?�4��?���}i�?�8@�@�?�{�'�E�?"�H� ��?Bc	2��? ��%iE�?j��d��?_Z�u���?�����?�"� ���?�y,Nk��?4ۼ�b�?��G����?�f\���?a ���?�qmL���?������?��� �?�e�w8�?�0��!�?@�8��F�?0��{��?�
�"{��?H�h%�?Tf��[j�?��D�#�?ڮM����?=�@(�?�J9;.D�?��k��P�?��خ"�?<V��'�?�肋�*�?<C�?a.��͍�?�y��b�?�Ѯ4X`�?C��%�?�hK|��?� x�)�??Q��G�?��(t(�?jK���,�?�O���?�Dڛ��? �:~���?؝�)���?Y9w�*�?�w���?V������?�j��@�?E�=��?���W���?l��Q��?߿�l���?5�"�?(:��/�?�zn�_�?z�W��?z$F��?��籂�?e\8���?NZ,�r��?�;��{��?������?�>�5��?�;^Z�.�?*QΗ�?���+
�?������?�=Ծ�b�?74�����?�Gے���?�'��R"�?%!��>@�?��+��?��LY��?�sh/z�?����Q�?��yQ�$�?{u� �?�����?Z��>Fi�?����^�?~=�s���?K��� �? +B!��?#�ڧ��?��傻q�?'(��l�?�=Џ��?�R��$�?"B���?�n�� ��?X���_K�?�$�@%3�?o�ۮ.�?Gd0cI �?:����?wv+S��?"wC0k�?�����?���%k��?n�E��m�?�T�f0_�?��\�G�?��"��?��ކ���?��2ui��?�-8+�?$ g ���?L�4�p��?� ʃ�?��V�V��?���>�\�?c\�ǋ�?���Q!�?\\�����?��@���?���O�?�XP�?�?������?����5C�?��#�Ѹ�?C�R����?Cw�����?�˴I��?����t�?��ed&��?�T|�m��?��j�;�?�҂`��?�4��?n���X<�?��k�ar@�����?w�i���?�FK@r�?D�,H�?���)I��?_�+G���? .h��?05;y�?]����?�A�9��?J�ɡ���?�!�8���?i���u��?a�sGRe�?q�����?��~ڝ<�?������?q�/��?E���?�"F�X�?�*���?e���?�؛0��?�����?۫�s�~�?�i>���?�-g$�?�\U����?"�NX���?{;$u���?4�p��?�!n����?�[���?�N�9[�?qt�����?��T�r|@�1K4�O�?�<�e�/�?#�6��?q����?�t����?���k#@�"�xH�?|i�?ˎF���?HH���?ٙ���?�pd�@b܆�sO�?	`@�X��?Ď�H��?���:x��?��4r�?�5���
@Mh��W�?�٣s�?�������?����
�?k5]��?����e@�k���`�?�{h��7�?�*;)��?#�b@L�?��^��2�?	��q@�A��?��@��?��:�~�?���2�?��!��?��A�@�v��s9�?P�A�x�?8�%K4�?��O_��?����!��?���ȩ��?^�wzp�?�I�)�[�?����?a|]��L�?���aC��?��-�P�?w��4�s�?<k=��?��9��?2�Z��?���pZ��?��o�!~�?�-c�?�bx,�?�,=�*�?��X�]Q�?�0�C��?��t�2<�?7m�!WQ�?e.�uY�?�o�����?����Y�?�~�����?��� �]�?w[x�3s�?���^��?_�ŘW
�?� ~F�9�?�ݺ����?!Jj���?V��9qv�?V���K!�?���p���?f��c��?�u�c��?#��K� �?�m{�O�?��\X:e�?�R�<=�?�P�cN�?�/�#��?���� �?Q5�ʎ�?A|@
g�?�+���e�?#����o�?� ̤���?K&>��?��&?��?z��xNi�?K�H| �?0�;@�?>�mw��?}��2ʫ�?��L���?���W�3�?[0�(��?a����?�a)�.��?�aJ'�q�?��L-��?L'&�x��?����E�?X$��I��?�a
���?����|3�?��q啷�?���~��?�����?�1�����?u_���?4�����?�?�	}�?�ÍS}�?�~� ���?�ބ��?z]�iU�?'�eJ)H@L�!�+�?o��?2��K.6�?���#���?~�?��?��N�@�}�[�-�?z�6���?�7R)o�?L#B��>�?�٧O�I�?V�r�e@ep���2�?���q�?�Y'G*�?�Nh߲�?P�H�)�?6m��\�@�����?l��^Wy�?��1bv��?ADu���?�J:m/�?xP::/�?L� q�?Xu����?B�}QL�?I��kȊ�?���11�?)�K��?��Vy�?U�i�/�?�8���n�?2i�;���?�U3�(j�? ����@�c,U�?�KFo��?���b*�?-�-NӤ�?�a�G3�?���qc� @�2�L��?��J�D��?�	���?��d���?�'/ǁ?�?�"� @�A����?�(��y�?0ݤ�	G�?�����?�F(�P��?�|�-��?*��ʔ�?U�"�/�?�#vߐ�?�c�,P�?����?�RS����?o��uL	�?Je=~
�?@���?H���D�?�"����?��}�� �?ɓ����?��M���?;���?�W��S�?ت֥_��?v�b��?N�7O�?���i]�?'�����?�ɣ/��?�k[��?�Ԯ�z@�71�e�?L
�Rs^�?�0�g8(�?�`p�o�?\�}	{�?�a�E�f�?CJ"�-��?�n�Ȏ�?�ܯh�?xB9?�>�?$|���?i]�RP@��A\�?�s����?RFH�l��?Լ%�?�)\3��?r���+1 @�t�;��?�ȚPL��?�9�û�?�j��?lnk���?�p�Kj2 @?��Ƙ��?�}�b�
�?�����:�?�i�o��?�tӇ� �?|�w���?������?<dݡ�r�?t�Ǳ9�?�V� �?�Ӽ��?J]�^*u�?��A�u�?����I�?��/Т�?¸�����?��%�j�?��p���?R���y�?/W�����?͈�G��?��r�J�?��Y��?�r%���?U��GN��?ب6�U-�?FV㕧\�?�\�$��?$#(ę��?���M%�?��z�҅�?�pݧ��?�C����?41y��-�?47���?�
}sw��?��Uۃ�?�;�K=��?�Y��`��?HEEY�?���<���?��ň�?_�L��?z/�V���?m��� @�����?$�aX��?6L�]w��?�O�Av��?a�S5��?j���7@<S��<�?��3w�?��2M�g�?���K���?\.�0�?�?1d�@����P�?�����?��mH�V�?�|��]�?�����#�?h$zɱ@�鑭Y�?/�G"��?����	�?����^��?���0�S�?Z�u��S�?}L�i?�?�"�c7��?^滆Rc�?�2����?�*���?Lͪ�W=�?I˺��?�;����?�s��k��?�c�/��?7bD����?��8���?6	w��?9�����?�ϐ҅�?�v�A��?�`��?�>
�2�?��N���?��6�ց�?�h]����?繩[*m�?�����?��T���?���x�?����"�?UKC�{�@<W�w&�?t�ݕ;H�?K��{j��?�q��6"�?�{mJ�?nNڗ�@��g���?�|٢@�?f�k�?h���@�?��{t*�?5���@\Y�*�?[��tC-�?�B��VX�?��>:�?�ؾ��;�?C�Pj�V@��~W�?�z����?�4�f�?�Uؗ�D�?��_����?!���9�?5I_��w�?�,ގX	�?����2��?%8��|�?�~AK�s�?Vfz��%�?з�a���?����h�?F�zH�
�?��%%��?å�z��?�V�1��?H��Px�?���(�?;�����?���B�5�?:���k�?��&�?j����?�s�K��?��v5��?B@:�WO�?�����?@]Гl��?�t/stt�?E֠��S�?;E�#��?]%�%�?��B�}�?�h?���?i�oۢ�?�uO�v�?H��y���?�0h�`��?;C�q��?3|`!Z��?�<����?\��Y7��?��΅T�?���O�?��}R�?5�`��,�?Q�~�?j�A���?11�PY�?�To_�a�?��~,�?��؎ �?��O�z0�?Keb�?.���.�?�����p�?C��b �?�
�|}�?7D�/b�?~w[�w��?�c�u{m�?rG�&�$�?A�����?h��ep��?��(�6��?�R�5 ��?��[rV�?v�ϗ2�?�a��?�ψeĴ�?�1^�	�?6�Z��(�?���[+#�?�3eW��?&c���%�?a��l�?�2��p��?G)JF��?��Ô��?��to��?3�5~��?�˃�x�?n�o$t�?�u0��?dO��?���?�Xf���?E�T��u�?+,�hw�?u��y�?$��5���?vC�1���?`s����?>�9��o�?I<���}�?V]�P�?�m8�H�?��`�sz�?qDtqEbX
   _n_supportqFhhK �qGh�qHRqI(KK�qJh;�C'  &  qKtqLbX
   dual_coef_qMhhK �qNh�qORqP(KKMM�qQh#�Bh       @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @�����צ�w�     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��ꢔs�r{�     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��9D����y�     @��     @��     @��     @��     @��     @��     @��     @��     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@��*E�p@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@k市�H�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@qRtqSbX
   intercept_qThhK �qUh�qVRqW(KK�qXh#�C�i����qYtqZbX   _probAq[hhK �q\h�q]Rq^(KK �q_h#�C q`tqabX   _probBqbhhK �qch�qdRqe(KK �qfh#�h`tqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh#�C�i����?qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKMM�qvh#�Bh       @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@���צ�w@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@ꢔs�r{@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@9D����y@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @����*E�p�     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��k市�H��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��qwtqxbX   _sklearn_versionqyX   0.23.1qzub.