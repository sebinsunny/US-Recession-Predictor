�csklearn.svm._classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX
   break_tiesq�X   kernelqX   rbfqX   degreeqKX   gammaq	G?PbM���X   coef0q
G        X   tolqG?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqNX   verboseq�X   max_iterqJ����X   random_stateqKXX   _sparseq�X   n_features_in_qKX   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
q X   f8q!K K�q"Rq#(KX   <q$NNNJ����J����K tq%b�C      �?      �?q&tq'bX   classes_q(hhK �q)h�q*Rq+(KK�q,h X   i8q-K K�q.Rq/(Kh$NNNJ����J����K tq0b�C               q1tq2bX   _gammaq3G?PbM���X   support_q4hhK �q5h�q6Rq7(KM��q8h X   i4q9K K�q:Rq;(Kh$NNNJ����J����K tq<b�BT  	                           !   &   *   +   .   /   1   2   5   6   7   9   <   >   ?   C   G   I   J   K   L   M   P   Q   R   S   U   Z   [   _   `   c   g   h   j   n   o   q   u   w   x   y   z      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                   $  &  ,  .  0  1  2  3  6  7  <  >  ?  @  F  I  K  L  O  U  Z  [  ^  `  c  d  e  g  n  q  u  v  |    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                               %  '  (  -  /  0  3  4  5  7  9  ;  >  @  B  C  E  G  J  N  R  S  U  V  W  Z                8   Y   �   �   �   �   �   �   �   �   �          #  -  :  ;  A  S  T  j  �  �  �  �  �  �  �      ,  F  [  \  ]  ^  _  `  a  e  f  g  h  k  l  m  n  o  p  q  r  z  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                     !  #  %  &  /  0  1  2  3  4  5  6  7  8  9  :  ;  <  ?  @  A  B  C  D  F  G  H  I  J  K  L  M  N  O  P  Q  R  S  T  V  W  X  Y  Z  [  e  f  g  h  i  j  l  v  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                 q=tq>bX   support_vectors_q?hhK �q@h�qARqB(KM�K�qCh#�B�W  Λ��e.�?�{a���?�D1[�U�?Z��Y���?�z�G�@��V��M�?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ��Ҋ��?
��Y0�?�G*;�?      �?������?��Q��?�-�����?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?�!ފ�?c����?��J%%�?��(\���?�G�z�?�~���?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?עWG�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?�*�N��?
ףp=
�?_�6�?:����R�?�p=
ף@}�"�>�?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?�a+� �?O9:����?�f^w�O�?y��x���?أp=
��?R��i��?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��K�?�&�j��?7��P^C�?F�����?q=
ףp�?��G�z�?:�5+�?��sr��?��3���?�V��?��~5&�? ףp=
׿�{�j8�?�X�y"��?%'¸Lr�?c�/�]�?,mG8��?�G�z��?�^���?�3��j5�?l�O����?�4`Zz�?n�s�p5�?H�z�G�?5�H���?Un����?�������?#�R���?]�����?�Q������j;����?���@���?��a��z�?�����?�5�3z�?H�z�G@������?!ml���?�9�n��?Ѕ�	���?��'q��?�p=
�ӿ�}G�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?�Fm�}�?�/Rm���?q�Q>	�?ݫ`���?=
ףp=@�+H���?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?\	# ���?�߈��?Ľ9�X�?и[���?\���(\�?b�����?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?ű�r��?�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�5�����?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�!�/�?P@��}�?��k���?      �?�J���?�������?"t�I�+�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?����?��R�y�?�����?�s@ڦ�?�p=
ף�?7���M�?�\7z�?���"��?����}�?7�j�?H�z�G@�N���K�?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?��O�V�?�m�02��?;r����?���	���?����<�?��(\���?�ca�M��?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,�����?�h��g��?O ���E�?��mQx��?��vY��?���(\��?`���+��?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?[�>���?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@c-�Gb�?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?v�����?t}ja>o�?\�-�=�?�Jpv��?��|j��?�������~���-�?���#�?��qPt�?���J��?�T�w��?�Q���?J������?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�����?^���*�?Z5�Uc[�?���l��?Ҏ#��?�Q���?��.?�9�?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿR��-�?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?��.����?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?c�2��8�?l�l��?�����?T��S���?�p=
ף�? ���P��?��H��?�z�G�?G��ֳ�?
݋н�?R���Q@X�C���?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?t��Y��?��1���?wF]�K��?={��?������?�Q����?�K��?<�	��-�?�U'�*6�?4�(�e�?�>���?֣p=
�	@|`�"���?�D̥�
�?�Zk����?��iz�?���\��?��Q���?��е:�?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@j��!��?�t&����?��(��(�?�^mSz��?g�Bg�B�?������@�5cJ�,�?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?      �?"&�H
�?�?�4��yO�?��)��?
ףp=
�?�=4Q�S�?�aݚ
�?(������?� R�M�?��7��M�?       @St��i��?���e��?I��/�?i�(�U�?�VC��?T���Q�?�74��q�?��O�?�\��\��?��_[�?fC�V�?���Q�@��8܅�?}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@�y��L(�?փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?����y�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�Ǔ���?ƪ+�K�?~r!�f�?�`(vo��?l��';�?�������? !�!���?�Ĭ~��?��Q���?>s=��^�?�����?�(\����?�a��~�??d~-��?�u�����?����2�?� ?7��?      �?��Ld��?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?ѳ!s��?�2�j���?     �?u�;�F�?�$I�$I�?�z�G��?Ud���|�?���[�?����NB�?b%c�r�?����]�?hfffff@Wd���'�?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�\��f��?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?�qV��?�z�G��?�	ϻ���?J��I���?�G�z @��w��?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?�h�(���?����?�3��=�?g�=���?�������?���w ��?Eb���?��Y@�H�?�|��X.�?�������?��Q��	@�ڱ���?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?���+*�?�-шs��?���ҋ�?�#o��?q=
ףp@N�Π21�?�}�!���?��Sڃ�?xE.�;	�?��}A�?��Q�@�=k,�y�?Шx�?jF���?������?�.�?��?�z�G��?��2}��?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ʞ2����?��	��?�jL�*�?�\�K	)�?U��t>�?�������?�ϗg�?�y]>d�?g;>)7�?�Ǭ�NR�?&H-/|�?=
ףp=
@VS�w �?�
�����?���!y�?��S��?�����?������ܿ����c��?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?6K�b0�?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?9�IA�?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@�����?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?x����v�?4H�4H��?�)~�r��?���Kh�?�p=
ףп�����c�?�$�l���?d!Y�B�?k���?"�?d�*|��? ףp=
׿F�w�M�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?�����?IM0��>�?��I��?�h�k��? R���ѿ��B+���?�v���?U�����?����?�M����?�(\����?2�g2��?�=�,;��?!G%޸��?������?ُ�؏��?�G�z�@������?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?�-{X�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�Y��.�?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ�5N�m<�?Za�T�
�?�1���N�?D��car�?�MҷV��?H�z�G@Ƨ�/5��?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?�_{��\�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?e�Y���?(������?�[����?������?��Q���?{�Z�˹�?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?�������?�m����?G��|���?E4Z����?�z�G��?hE�-\�?
��\���?��\AL��?)us�?      �?433333�?@�����?�e�:�	�?Dy�5��?��:cc�?�b�X,�?
ףp=
@�j��s��?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?���p9�?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?��9k��?��i�,�?ףp=
��?���b��?,Fڱ�?��Q�@9��V���?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?�~�A
�?��0��?R�}�=�?ӗYl�n�?.�袋.�?�Q���@N��i�?s��&�?(W�7�?���xW�?B�HV��?��(\���?�LGuk�?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?կ~_�:�?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�?뚖f�?1ܫ`���?��Z(~�?�;�;�?@\���(̿O�e���?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@C���P�?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?"K�_y�?���,d�?���<�?jhɬ�?�Q���?D�&Dq�?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?����S�?�N�u.�?�&$a��?���7�?      @6�� ��?W����?��8��8�?      �?Au���?�������?(Bo*��?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���? �X��?
ףp=
�?�Ѣ�ǃ�?�;⎸#�?      @3����?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?'���/��?��
�	�?:[���:�?�!!?�Z�?�0݂k��?�p=
ף�?̓�lXD�?{���T�?=]�΁A�?�DJ#��?���e�?|�G�z@��F �?ϙΔ�?a#@i��?M��d�?��,��?      �?;���?�wF�?��D'�?6������?�_�_�?�������?�Ko��?I��q��?�'iq��?�&��?#�����?�Q����?�E��Q�?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?K]E!�6�?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?����g�?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�vף]��?��;�l�?��{����?��`|��?���!�?@\���(̿Z�S�Ҳ�?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?PPvI�?]�����?ea����?m۶m۶�?
ףp=
@���UY:�?��Lf�@�?�!��uy�?������?�aS���?�G�z@���{��?�p�|���?���)��?^�3���?h�J� :�?�Q����?���ah��?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@��j>��?��+���?G]t�E�?X?A�x�?Ӱ�,O"�?�z�G�@����� �?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ(�~��?�>����?      �?0`z��Q�?'u_�?�p=
ף�?W�n��~�?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?�a��P�?��#�N�?{�G�z�?�A+珽�?���9��?\���(\@1O�u�?�N"H��?����?Hx`2��?��r:���?������@�P	�_�?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?�����?�Qf�,�?z�<���?�%���x�?Z���(\@��w]�f�?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?vP�I��?E8S8B�?������?�5��P^�?����������(�?��I��?      �?	)�L��?ڟ�!T�?��G�z����8I;�?}9�ot��?d����.�?֐��<�?OP�?�z�G��?�dn�>�?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?/G�9�?�����T�?`�t����?	�m?���?��Q�@�J��}��?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?�܎h�?��/�$�?�p\��?���6�?���(\��?�=
��y�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?�j�с�?�dn}�?�xJ�Rn�?��寖�?�z�G�@�s׾�?:�SR�?���7���??	-zռ�?��y�?�������V�o@��?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�w�x@�?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�?��*@�?:��8���?�O�Xs-�?���#B�?��Q���?��;���?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?:��]��?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?P�ϸ=�?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?�83���?�{Nm{�?�F�� �?�������?P���Q�?1l(�?erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?�J/��?e�F-��?�������?���:%�?V���g�?ףp=
�?´�z�)�?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?2�7���?���A�?���i���?_7��T�?R���Q@yJA���?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?x��l��?Ɏ �U�?�˴�`��?��N��?`���Qؿ�zz����?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?�y�]��?]�)~I��?��@��[�?�{����?���(\�@#i��K�?"�FU��?�71}�?v��3���?�N�Q�S�?�Q����?�5�,[�?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��A��?�P�6Ԗ�?s>�cp�?�`κ��?���$D�?P���Q�?爈��P�?���\�?�^o�?�?Q�/��?^̧^̧�?�(\����?�XrYǾ�?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?�X��e�?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?J��YL�?VUUUUU�?!��a���?�7�7�7�?      @%CE����?V�gb�?��W�l��?U�����?_�HI��?�������?��h~3�?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�<��2��?ӏK�K�?��{���?���S��?{���g�?P���Q�?�Z(O,k�?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?�
>U�?
ŭP�
�?Pf�i���? i]���?�G�z��?�_����?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?2E�Ĵ�?	��-��?'m�`�?:o1���?hfffff�?��E T�?��j�G�?u�5�o��?���d��?�~��?�G�z��?\�o�nl�?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?��mW(��?333333�?"�*|��?���?333333@��K���?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?�צ����?3�*�" @�#�p�j�?V�;^l	�?(\���(��9���r`�?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�	ږ@��?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?��h�D��?��P��9�?�1$0��?}��O���?833333�?&~��.w�?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�s����?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?�o��5�?O�o���?�7��ֲ�?J"���?�(\���@������?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��??V�)��?_�_��?      �?��B�
�?�G�z�?�Z�K9��?�SR�&�?}�K`]�?��<d��?w�C�v�?���Q�ο�*UۄP�?������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z���c���?_������?���h��?�����?\t�E]�?�������?LkCJ[�?^e�NF��?�}�K�`�?GT��a�?&Դ���?P���(\�?iS�}s��?KY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(�w�cK��?�q� .�?��"E��?�V���2�?�^�^�?�G�z�?Hݽr�?��]���?[�[�@�{�q�?.q����?���Q��?�@����?gDAl���?<e�U!�?��-��?'u_[�?�Q����?"�R[WD�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�?�S�����?���NV��?��=��?^���?��Q�@�D�y*��?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?�Gq���?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�6jDRf7�? ��2�?S�n0�?���&�_�?I%�e��?�������?����5�?w��{���?)�b���?z9��E�?�0��=)�?�������b��i"�?�'���?�*H^�?�����?Oozӛ��?,\���(�?��x~q��?�G����?h�[�t�?`o�3���?C�l����?
ףp=
@�T��T��?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?y��RE�?n,�Ra�?�$\Z�?��S�p�?�������?��p�4[�?T�.�n��?�-�׮�?H{����?������?P���Q�?��/>�?Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿ���?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?���6���?�w���?zkfkl��?�k(���?      @�q�^��?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�X�!)b�?錞�m��?uh���?���g{�?���5Q�?P �9� �?W�4�d)�?��AA]��?�E�)}��?D0���?�����?%'#g��?�Q��?w}uUU��?b���?6���@�?��e��?����_��?d�F
%�?}����?({{����?N'�܀�?�X�[2�?V�8"}��?�t5�^ �?f�w��r�?gsT� ��?�7}M/�?Ո����?qM��=��?Z��OY��?����Z�?�0��4�?5Z��D�?�,3�&C�?�h�Ѕ�?Ĺj���?\�ڈ��?\��>�?��G���?��mG�?�����?ݯE��+�?�|��U!�?��믽�?}wQN�?l�r$��?���I'��?�ѪCe��?���p��?�]D�(�?��6�}�?�� /�?E�O��?`�B��?4��+,�?�ӑ6�m�?o��ߝ�?�=	p@Q�?xE;J|�?b��"�?T�T��?ʹC�H��?����;�?&�x�|�?�g�3S�?��E&l��?q5=���?��[�)��?��	���?�Jx�4{�?yO)+���?�m�� �?-��i��?/i�:~�?Li�ǽ��?�5rD��?*�(I��?  �F�?ٌ�
���?��Fy���?�Q�?��Fl^�?��� ���?�����?8��Q���?L����?�_����?��^���?�tX��?"h'j9�?�yڿ���?��z�6�?�����?�P��	��?����?���*���?+�Q_���?RcM[T8�?nK����?�_��	��?e8��+��?k�L�%��?y �n��?r9��-_�?�H�v��?�~�M�?�!��5�?@�JmU�?�P�d��?�:�(��?(��	i��?�-FO(��?����)�?FQq�EJ�?���*� �?�%���#�?�9�����?3	��P�?9Ʉ7���?!s�`S�?��j��$�?����-�?�!g���?�V�`���?�ƒ�/@��YoZ�?B{}�N�?eR��ް�?'̑[�!�?a�U����?�R��p9@������?���]���?���\�&�?��/���?��|M��?_��kB@������?uF6OeV�?0��8�s�?W8}��?���<�k�?r=#@b������?�B�2��?WL�1�??r#���?���{B%�?V�v�p@U9 ��?xp�0Q�?��&,��?}�� ��?���+��? �VR�,@>w���?U0m�<�?²���?��j����?,��9
�?��A1@�z*���?�	�v��?\n����?��QJ��?�.�?�̫)`@�`�L���?3u���l�?&B�+:��?�����?�d�j�?�V �@$G�s7�?{D�^��?nf���n�?=���m�?O�x$P��?x�m�E��?�W�[{�?�K �?>S����?��ل
3�?��y���?	`J��?}ׂȑ	�?�8��N�?�����?Q{o��e�?�>�:�?Q㜷��?#���?8�Ow��?�=����?F�ZK��?�9x�?+V�^�@�o�S���?{u��2��?%�����?J2�5��?�TÑv7�?��CK@�ا�6��?h��;`E�?�����?��N����?n<� 0�?��uJ&@�k�/ �?,�u�UF�?��	�?�AT.�?�q����?��/�@5� ����? ��XMn�?��Tt�O�?O_K��)�?5^8���?��:d�@7�u�fX�?�L"��7�?�'�S�x�?U�6��?{)AX%�?���H��@q9�N��?�]j�;�?�lw�Bl�?z=���?V�L���??���H@�������?־���X�?�3�����?��_I(��?�D?��!�?�6?r|�@���mE;�?�Y�=�?����?F�oejl�?��F�M�?��5ǋt�?�!�%�?Rh��(�?�����?��$���?%�!���? �˝Z�?8܅Y�?��݊���?�B\~g%�?���H#�?u��,�?�5Q���?~-�<�?!��R\�?L?�<A�?\-c�?��@c08�? ���Yu�?���r�	�?���sT�?���/��?na�y|�?G�Ɏ(�?�W�Ę�?���R���?z�x�?�"�c�?M�E0E:�?6��?�(�^���?i���>#�?��V�g�?ݵ����?p{��g�?~���?��{�if�? ��,X��?M���l�?2����;�?L�➖7�?�
��?`a��˼�?�l	#���?��s�dR�?R+&����?�J
�I��?ݍc�-�?] ���K@x7��>��?)�v�?�?������?�@�?�?I���T>�?�߅���@	�V�D��?*�B�>�?�^D� ��?�p'
�?)��O��?z9�f8�@w��<.�?�ayqi �?��[���?3 ��)��?vdS}�?�N�K@�%%_�j�?�c�9�?��qP�?2!E=���? �`$*�?�fuG:�@w�W��?�@}��!�?p;���?�.@{���?�+�d��?͈��p@Pwd6e�?���,'��?��HJ��?^�8���?0�����?��ܙd*@|j(���?(rت&�?/Gx.�,�?)�ΐ���?�����?�v3�:@�����S�?z��IT	�? zK��?~���O�?���Z���?�h�x�N�?�u����?����{T�?�.��8�?�d�aP�?ހ����?����H��?^$����?�x�8^^�?</A��?��x��?ל�|��?�9g*�>�?�kg����?� �zT�?e��q_8�?NV�_P�?%�V���?u��A���?���o���?cqN�]�?>�6n�?�"��?ݼ�܀C�?@l�xT�?���2.��?6��M��?LX��~6�?�����?�c�����?0�a����?����b�?�*�r^�?�E��?N���?��T���?����P:�?�|#��?'�0��H�?>�xK��?�9$l�?��u�o�?�Mh\�?�Ŋ�m��?Wd(�T �?�, ����?WPw��?�l/�?���>���?F�`؜��?^����?�(w���?=~�p�?����.�?��P�
�?H�%�e��?��I y��?��x��?����0��?�蠶wE�?�x�.���?��d��/�?J�p%�?���G�?�V^�z�?4M:�?�?>�7��Z�?����h�?X�����?k@���R�?����t�?�̤~i��?��s�(�?�����?fe����?=#�f�?���@�[�?�d�����?�9�;��?$v����?���R
�?0�J��l�?9������?zx�s�?a���8�?Ւb����?���z(�?@�9G���?1_� !��?��?z���?;������?���=G�?~F䚰��?�%���J�?�YX�m�?l
WjCQ�?���)[7�?�oqe��?��H��?g�	�?����?�;=��:�?�zS1���?ڝnm��?�\x�#�?(�wydU�?H�UM�?A��ܹ��?��x<}v�?G�����?�%���/�?z�޾�6�?�
�p\�?��벢�?��/���?��۪�D�?cE�LK��?n*�F:�?�Z�*�?3eb�?'Ĥƈ��?z�� F��?b'R�^��?]�ި�?W���"�?�p�r#X�?���Z�?�(&�K��?����#�?㢓�rU�?/�s�NM�?�������?�E�\v�?{�,��?d��q�?U��W�?x�*�݈�?r��?�P�>{��l2��|�?	_6#�?AHj�h��?��L���?͹��a%�?GR�Q7ǿ(oi�a��?C�����?��ŋ��?�2$�	�?�_��k�?бc	�ӿ�� ���?�]fs��?��W�?fӺ ��?���S��?l���տ��1�?���L�?��J,Ӝ�?�}��?�?9~?���?.�O��M��O��^��?��,��?�*����?8���?牑�_��?69���?�/�b,��?�_e(�?C����?S���7�?�[��S��?�ɾ�
�ҿ	�����?X	���?*�M�w�?�_�jT�?��:�u)�?Dk���}��+:ٷe�?4׬[��?�ƌ��?���%��?�4"��o�?�ygX(+ĿA)�[�a�?.wO��?k 0u�?�~��ǋ�?�2E�]��?�1m�#���ĹM��?��D ���?�H��s��?P U�7��?���N�?��e Rſ�M�g�M�?���bE%�?h��|�?�tCӪ�?��a��?Ik���˿�{�x.�?���I��?	B����?-_�-�?��/�&�?K����?�U�3�6�?� 	g���?�t�B/��?`�^��?&ȥ�|��?�G���8�?�g��i�?��[�=�?i����� @uS�j���?6ST�*��?̠��E��?��&��O�?��V�Ͽ�?4
�>�?�m�tU�?rNx|��?�����?�M����?��V��G�?��-�ԯ�?�#e-�?�E�/�#�?<���e8�?B�h���?֥*f ��?;p��N��?�^O��3�?���#'�?�T�#��?3J�P�^�?ז�1�A�?K�yy�?�����b�?�ϩ�)d�?`�[����?<�J�?�4|@�?=�r�o�?n�*���?���U`	�?\e���r�?j�����?r�����?\��?Y�2)��?Ιj�x�?�Zz�~�?Sl�W:Z�?nGa�!�?�w=���?�>�� �?� w2�~�??��qg��?��|'pg�?���/.��?�9�s @�v�æ��?�f�7Ɣ�?��z����?������?A�*b_"�?�_4�U�?��ۘ4�?����\�?�<0s��?��;]��?0��9��?��uǯ@j���q�?���9��?��`eq��?�a�Jr��?��	�RN�?�慍N�?���Q��?1��?GcA����?P�!mZ�?����s�?$��$�?ݱJC�?,z]t3�?m(��4G�?���!�S�?� �����?���`��?��a���?~]3ne�?(��>@�?�7��t�?e5s�W��?���m�?�2���_�?���e[�?�SA���?��D'�|�?�4㩄v�?h �ƭ� @'��T���?�Z-i���?�y�JE��?+�C˧�?��n���?�쥡��?����h�?{i�c89�?! Rf�?)��W���?*���� �?e9����?Ҳ�U7�?�,��K�?5�a秶�?+sD�ѭ�?�:�� ��?��L����?�T<�׊�?��_fߐ�?F�!Kd\�?yZW��?����Q�?1&HZB�?()z��>�?q�GZ�$�?�[.�غ�?7�M ���?��Գ�?. ���?\;I|�?�� ɸ�?�l_f���?A�%~vR�?���4��?);�*��?��z����?#���?-�J,@�?����O�?�4���?�l�s��?�ͩ�ܘ�?�I����?a^�|��?������?*�5�R��?m��Q���?ׂ����?dz���o�?����H��?���}T��?��D�V��?���.�r�?�hϿix�?��'��?�w��?��پ��?��0�jL�?T�H@���?s�}F�c�?��&�?��8X���?�X�Z�?=�G]�?��OK<��?��X�4�?4����?'ޡȧ�?������?�;�,9s�?�(B�>��?��STu�?���5���?����g��?�Ր����?_$�-���?��6}a�?Na�d.�?��b{8�?�2�ɩ&�? �f|�?���ת�?`��jN�?Q+�-�?`�:��C�?^�͢��?/�!��?x����-�?bm�Z���?vc��H�?B���h0�?f:�߭�?��;���?������?	�[�k�?�v�I��?�:��޵�?-�\���@:i��a��?Ŵ�'_��?��:?��?TJ�ok�?�M�;��?(��{�\@&�2�D��?�[W�֘�?����V�?m�C?���?�DA1@L�?IA�hH�@���S�?Q�3�y��?l�Fp#��?��p�h\�?�?��?�S��NX@<��h^��?�w��O��?��C����?�����w�?�Ԑ���?�Y�ײ@;}��]��?�➯
��?6 >v�?�a�����?�=��6��?���'@\g��N��?R�{~��?(d�����?������?�BCӧa�?(qoO�@�Տ�6�?Z\�3�^�?~�Yn�?a�FNT��?�.{z?�?
ܵ��@��&?z��?�
�-t��?,s�
`��?ޒ����?����w��?=?���E@~,o8���?��$Y���?)�t��?���5���?�< ��R�?F�B8�@G̻��?�ܮ�Һ�?%��[�u�?GAX��w�?$,�b0��?�����A�?G���%��?��*����?SSqC���?��H�o��?q��n�?Y��R��?H� ��? ����?mr��w�??�2�x�?#E2���?����:�?c�ap��?�б��?Wܲ��p�?�⅌X�?~|y�0�?1 '���?V*u��?�Cq����?/B��g��?�^����?�1l�O�?N�w���?c~��!��?��E����?�n�&!��?=0Z�|�?�M����?f��lK��?�>e/��?����^f�?0c��*��?��W��g�?��o�G�?��Қ���?���t�?S��s&�?���v>t�?��]5�?0x�$�=�?	 �	X�?OE�yj��?*�}X���?�Yº	�?�?��E,�?�kO����?�~ִl��?���,} �?������?J������?A ���x�?����'Z�?�p�!�?��ɾ.��?�ܭ\6�?�@���?n�{�?�?�0/,�?:Q�+���?��(1g��?�Sür�?(N�9��?�v�t�?�������?��{�k��?�ǉW��?�V!�I��?�̇����?أ��>�?�\s>#�?]����?�L8�4�?x�����?�H�V(;�?Q�����?���Q���?G�.}��?�6���?�@8�"�?)~-T!��?�e�a�?~�-��?�c��6�?ª�����?�}�b �?D,�p��?�{i]�!�?�Y�.���?��,�Q�?�l8(U�?
��$��?w2s�G��?`�1�v�?�`�v��?�=9��?��n���?Z������?�UR����?�a�W��?��)����?�������?)�����?��!y9
�?�m�]*��?��|8-�?zF�����?�]��t��?<VOԯ�?�Dw0@�?���]4��?h�^j�?�f^�5F�?�zR�I��?��z#�\�?������?��n���?��~J�?b�#\��?�{�d{s@�Ȁ࿶�?�rv	 :�?��]���?��?��?�;�Z���?b1���I@v�ɡ!��?��rze�?�A��'7�?���OE�?�?�W��?K����d@�P���]�?�Թ�C5�?� Q���?g�rO���?|]���?~M��
@jb"ʁ��?�C�<
��?+þ̜�?Z�@��?ִ�<���?�M�@&�@��'s#�?�Ao+�?FlN;;��?�?ے��?��b�z�?���nl@r/��-�?��E���?��/p��?,d�:	�?�y�_#�?s�)m�H�?���1�}�?�x���?EA|p��?0x����?N�;���?�F�T�r�?Ղv���?�߅g���?���㤍�?cB	Y���?by?�{j�?������? A�Z�?�d�A
�?�P�C`��?�$x��?l�
E)0�?��к��?_�#��?v(��'�?������?�$=��?� D��P�?��Sv��?t�fa���?��`����?i%����?�P�`���?�R��.�?5v��f��?���n��?�!��~��?����5��?��=\�?c�9/��?$�x���?��c�?��<"2��?L�?����?�6L���?�^�U^
�?����'�?ܔ+d�m�?o�(|�?$7e�7�?�x�a�\�?��qy_i�?��o��@շQ�?������?�?��d�?">0���?-��ή�?�@_I8@�0�֣��?Ҹ8l���?�>g���?_��$��?�v~pp�?ʶ[�L��?� 7Z���?�җea�?l�,�Q�?QųR+��?5�(�ſ�?�e�a���?��H!uP�?��]g:��?�IS%�7�?�O��O��?�;C�Y��?�AL��6�?Q9��?�Y2;Fw�?9�F/ ��?I �X(�?P����?����?��m_��?T����/�?�Ǿ|�T�?����$��?����?ޭ��Wa�?p�`���?\غ���?��� ���?y��}��?�q�����?��'U�K�?{�VU�?�6�����?܃��j��?Χ@����?P�:)�0�?�`����?�y�W ��?-0���?�X���?s(�����?'�����? <�r�@�?�˙�b�?��d
�?S$R�.F�?��0�D��?N����?�{���#�?� �])�?炎���?�]ښ&��?�s�j���?�����?��B���?��(��P�?�����?m�@�c$�?	GR/k��?d�8��?�vP����?B�Q<I�?���Y���?e��c+�?FN�/��?0��v��?��]��?����w[�?*OQjN��?�UL�P��?���o��?�ǀM�?���dɿl�$���?ט���?P��V�?&�*,[��?I[��Ch�?�m2v��?td.}�?���.��?�Ks�j�?Q�/���?qQ�d��?�
�Y�?K50���?��ۺ�?@ �����?�p�+S�?����7��?2����?�3����?q	��q��?GKEbN��?:�r�݋�?l��4��?G��m"z�?�4æ���?�_P@���?���'�?Ţ>x���?
�2n͍�?���50�?=��Y.�?_)�Xӿ�?�t���?���]�?iD�� ��?خ�
���?�P{�N#�?�!�lt�?9l�+��?vw�C(��?#��^��?x���n�?�:n�)�?�\��&��?�O��n��?*2�{)��?f�{Ӻ��?����!��?a�����?�l�+��?�-`���?�G����?9�&�j��?]�t�P�@�bR�?m�_I�|�?�շ�A[�?b��C���?
zb�̎�?ʛ{�b0@���?��?R�s���?�ާ�*�?�D�V��?���s�?�����?e��q�?sd���?vg;����?��2�/�?a쬤���?��N���?�qL�6��?.o'\��?tBW����?al���?��;��Y�?�!]���?����n��?�-�+��?+ת���?\��`��?��ni��?R.����?O6���?��>_"�?�O�޵�?�%:��!�?1�t}�?�=��y��?V�c}�g�?qDtqEbX
   _n_supportqFhhK �qGh�qHRqI(KK�qJh;�C�   �   qKtqLbX
   dual_coef_qMhhK �qNh�qORqP(KKM��qQh#�B�       @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @���-3�Bo7�     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��ΒF����     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@�x���{�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@m=�3�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@6}x�g�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@���!��V@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@qRtqSbX
   intercept_qThhK �qUh�qVRqW(KK�qXh#�C��
ѱ@�qYtqZbX   _probAq[hhK �q\h�q]Rq^(KK �q_h#�C q`tqabX   _probBqbhhK �qch�qdRqe(KK �qfh#�h`tqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh#�C��
ѱ@@qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM��qvh#�B�       @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@�-3�Bo7@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@ΒF���@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @�@     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @���x���{��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��m=�3��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��6}x�g��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @�����!��V�     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��     @��qwtqxbX   _sklearn_versionqyX   0.23.1qzub.