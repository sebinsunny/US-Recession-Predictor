�csklearn.svm._classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX
   break_tiesq�X   kernelqX   rbfqX   degreeqKX   gammaq	G?PbM���X   coef0q
G        X   tolqG?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   n_features_in_qKX   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�q cnumpy
dtype
q!X   f8q"K K�q#Rq$(KX   <q%NNNJ����J����K tq&b�C>���3�?���Ě�?q'tq(bX   classes_q)hhK �q*h�q+Rq,(KK�q-h!X   i8q.K K�q/Rq0(Kh%NNNJ����J����K tq1b�C               q2tq3bX   _gammaq4G?PbM���X   support_q5hhK �q6h�q7Rq8(KM�q9h!X   i4q:K K�q;Rq<(Kh%NNNJ����J����K tq=b�B                                                                     !   "   #   $   %   &   '   )   *   +   -   /   0   1   2   3   5   6   9   ;   =   >   @   B   D   F   G   H   I   J   K   L   N   Q   S   V   X   Z   [   \   _   `   c   d   e   g   i   j   k   l   o   p   q   r   s   t   u   v   w   x   y   {   |   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �               
                                    !  "  &  '  )  *  +  -  0  1  3  5  6  ;  <  =  ?  A  B  C  F  G  H  J  L  O  P  S  U  W  X  Y  [  ^  a  b  d  e  h  i  j  k  l  n  q  s  u  v  y  z  {  |  }    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                                   "  #  $  %  &  '  )  +  /  1  2  3  4  5  8  9  :  ;  <  >  ?  @  A  B  C  D  E  F  K  O  Q  R  S  U  V  W  X  Z      	      (   .   ?   A   R   n   �   �   �   �   �   �   �   �   �   �   �   �   �            $  %  8  9  K  Q  Z  ]  _  p  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �             !  0  G  H  J  M  T  [  \  ]  ^  `  a  b  c  d  e  f  g  h  i  k  n  o  p  q  r  s  t  u  v  w  {  |  }  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �          	                                         !  "  #  $  %  (  )  *  +  ,  -  .  /  0  1  2  3  4  5  6  7  8  9  :  ;  <  =  >  ?  @  A  B  C  D  E  F  G  I  L  M  N  O  P  Q  Y  Z  [  \  ]  ^  _  `  a  b  c  d  e  f  g  h  i  j  k  l  m  n  o  p  q  r  s  t  u  v  w  x  y  z  {  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                   	          q>tq?bX   support_vectors_q@hhK �qAh�qBRqC(KMK�qDh$�B��  �L���z�?X�O���?��F�{�?!���c��?�(\����?�g����?��=Qr�?7r#7r#�?y�sJiM�? ��c��?433333�?�Qa���?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?鄣Z��?:�SR�?���7���??	-zռ�?��y�?�������V�o@��?u�-BK�?��T��K�?��x���?>���~��?���Q��?f[t��?����?��Pp%��?kub�Q�?̟�Ѐ%�?���������X5�Q�?h�����?��1����?�IF��?�_{�e��?��G�zĿ� �����?{^Q�h�?       @��Tf,�?�7�7�?�G�z @'�oz��?��=�9�?�[��"e�?�+U��R�?�Gq�>�?��Q���?��� g�?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?��k�<��?�k��%�?^�4�y�?��xN%�?433333�?pjh����?��״��?Ѻ���@��O��?����T�?���(\��?���7 g�?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�?%���y��?a8B��?�!!?�Z�?���q6�?<
ףp=�?p�n=t�?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?g?�V.�?�aݚ
�?(������?� R�M�?��7��M�?       @St��i��?�S�����?8�P\�?��;^�?M�*g��?\���(\�?�	�;D�?\��Rx�?�ۚ��?�<�}C�?����C�?H�z�G@H������?yϠ�%�?      �?^���т�?      �?�G�z�@P��+��?�b�)U	�?�s���?�M�isT�?N1�^�?q=
ףp�?D����?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?0�|L��?�GZ<
�?�s�9��?�g�M���?���u;�?)\���(@����B�?i�+s�?333333�?`�>��R�?��.���?q=
ףp@=�f{?��?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�??[�w(�?��_O�?��G��=�?�!|����?L��7���?033333@�P�S���?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?*��Al��?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?[��`��?ك2�*j�?� �;��?�������?�(\����?,evp��?�@�,��?I�$I�$�?x�?q�?u<@�La�?\���(\�?�?i���?Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿ���?'�CU$
�?      �?�t�U�%�?.�#EC�?��Q�@)II��?���,��?ى�؉��?��� W��?{�G�z�?*\���(@�)R�?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?����=��?|�Zj�M�?������?���;��?�p=
ף�?��"�$��?Q�����?I�$I�$�?���Y�?z��!y�?333333�?ęmI�?�'=��?��fě�?��Xf[�?���¯��?�G�z @���#��?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?8K����?�9vZC��?X7�"�u�?A ��X�?ƃ'��?�G�z�@��n���?t��!���?,�X��?^*��U��?�:�>c�?��Q��@��K49�?���\�?�^o�?�?Q�/��?^̧^̧�?�(\����?�XrYǾ�?���. �?i�`���@jڪ���?��}ylE�?�(\����?ڔ��ɣ�?��Sr��?U����?<����?w�{��?<
ףp=�?�c��o�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�9��-c�?X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?��S���?V�gb�?��W�l��?U�����?_�HI��?�������?��h~3�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?F}�p �?������?N6����?\����?ffffff�?�T����?z&�����?�H(m���?��K�y�?���cY��?��Q���?��ʦ���?��B\&�?�n0E>��?���L�?2 K��?�(\����?O(���?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?�74J�_�?*6\u��?�$8����?�/t���?      @kp����?�!ފ�?c����?��J%%�?��(\���?�G�z�?�~���?)��h��?UUUUUU�?�����g�?�X>b��?���Q��?;w�9��?KY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(�w�cK��?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?��<���?      �?��(�r�?��a	G��?���(\�@n.>��	�?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?^e�NF��?�}�K�`�?GT��a�?&Դ���?P���(\�?iS�}s��?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?9�IA�?��Zb��?��+x���?� �Y]��?����?hfffff@N~��I�?�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?��m����?ӏK�K�?��{���?���S��?{���g�?P���Q�?�Z(O,k�?�4��
:�?(6$�)G�?(��J+z�?v��4��?���(\�@_�QU��?쟜�ث�?�$I�$I�?Q�d�?J��I���?0\���(�?4::RDA�?P,��v�?�������?4:�$�x�?�%����?�G�z�?Qj����?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@c-�Gb�?{��*W��?     @�E!��p�?�$I�$��?�G�z��?�_�����?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?P�ϸ=�?����8��?��*H�?>���h�?�؊���?$\���(�?X��WI�?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?���|7�?ۍ}��	�?>}���?��ũq�?��������?:��z�?���]�?��g����?1sJJ��?��f$/��?���Q�@�T��5�?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?�O�C���?y�5���?�V�ޑ_�?%���^B�?=
ףp=@�d:ޕ�?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?עWG�?m��C�?      �?2zW�]6�?��L��?���(\�@��y����?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?��L�F��?�Q���?6��<�?@(��?�;�;�?أp=
�@���d�?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?|? ��@�?gDAl���?<e�U!�?��-��?'u_[�?�Q����?"�R[WD�?L��,�(�?}�>C��?�t��l��?('����?)\���(@6J�!���?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�? �	�'��?pN�F��?�^mSz��?�]�P�?�(\���近x����?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?y���t��?a�B��?�������?' Z�u�?�����?���Q�@De�&���?�ӄ���?R���Q@���K���?����*��?�(\����?I^J��?����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?]T�%,u�?Ե7�rL�?�l��l��?���'��?��E���?��G�z��Ψ}Ri�?�o�����?��%�̀�?�\"�0�?P[AG:��?�(\����?*�(��?%n����?      �?7��S�?��/���?�p=
ף@�N�w��?"*����?�q�q�?�s�̫~�?+1��JL�?�p=
ף�?���U�g�?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?^` 5��?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?%����?��{�A�?,˲,˲@�Z�rf�?c��0u��?���Q��?��v��?�����?�MA�1�?I �����?,|L���?�(\��� @����?��L��?�q�q�?G`3�!�?O���t:�?R���Q@���Bco�?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?�צ����?3�*�" @�#�p�j�?V�;^l	�?(\���(��9���r`�?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z���c���?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?y��RE�?n,�Ra�?�$\Z�?��S�p�?�������?��p�4[�?8����?�gS��=�?�~��H�?�Vi�_�?�������?�11�G��?���g
�?&���^B@���X^�?��FS���?G�z�G�?;��q�?�_����?      @����,��?[�o�W��?���Q��?zI%D;��? �5�0��?�����?B �Gey�?r�q��?��Q���?���I���?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?�h�(���?����?�3��=�?g�=���?�������?���w ��?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?g�\���?�����?��񍔎�?����.��?�G�z�?'�����?�D̥�
�?�Zk����?��iz�?���\��?��Q���?��е:�?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?��m��?����?&z`�5�?2u�=�S�?      �?��]�E�?l,����?gH���?���2G�?v�A����?�z�G��?fÿ���?Jt_�h��?߈�N�@(���'<�?ZZZZZZ�?�G�z�?ۇ�����?��S3;��?ĸ_�T>�?��a8%��?�,�י��?q=
ףp@p��8�?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?���/�?�":>ɗ�?���ע�?���'-�?�R71�?      �	K�����?�n���?H���x�?6?�x�o�?�#�	<�?R���Q@4���'�?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��K�?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?Ŝ�lK�?."t��D�?]t�E�?N����Q�?�^�^�?|�G�z�?��w���?�v5C�?333333�?>FX�v��?$Zas ��?���Q��?�>��/��?n,���$�?����b)�?A�쎑��?@�1���?
ףp=
@,4�����?�#tT��?®b�?	�e^��?�m۶m�? ףp=
�?�)�9�?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�<��2��?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?It���?"K�_y�?���,d�?���<�?jhɬ�?�Q���?D�&Dq�?�,��o*�?���tT�?Eg���?�@i�
�?��������5H<^��?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?�-{X�?q����?*�3��?3iM��h�?QJ)��R�?=
ףp=�?��U#3��?��p����?      �?��e�N�?�������?R���Q@>����?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?�u����?�wK�?��?�ef���?tT����?�z�G��?��-��?�x�\�?��2����?ؔ�
&w�?      �?أp=
�@�t�#���?��B~���?ƶ#e��?-��k4�??&ǒ::�?{�G�z@8f?�?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�`1+�H�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?�d����?���-���?_l�9��?L��N���?P���Q�?�ON���?%��d B�?颋.���?N�|�?$I�$I��?�p=
ף@�3�V
�?=B�k��?g�K1_h�?;9�=-�?$�D"��?q=
ףp�?�D�o��?s����`�?�0�0�?��e�s��?���]�(�?�������?ApMrx(�?�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?#��3�U�?J��:���?=
ףp=@��=!E�?���E�?=
ףp=�?O����?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?����Z�?r��Z�@� ��r�?g��|�Q�?033333�. }0�b�?��TD��?x!�����?�x�;���?���&P��?�p=
ף@3�l��?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?'���/��?�'Z�:��?�|ۗ�s�?�#%Ŀ�?�J�gQ��?��(\��@��^1���?T-����?UUUUUU�?L�5���?�������?ffffff @Ι�p|�?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?����em�?׊��+��?Y�����?"$�A���?�(\���@K������?F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿr���;�?-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?�X��?w����?     �@R���8��?�~|���?P���Q��u�%ܚ�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?�՜�pH�?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?�X��e�?EÓ���?�����?�&z��V�?WUUUU��?���(\�@$i��!��?֊�q��?��Z��Z@�K��?#e�����?���Q��?
k#w��?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�	ږ@��?�r�4�?�;�;�?ڡf6�K�?�s�9��?�Q����?�+F�d��?���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�?�k�6��?���~�?9"�P9�?<O�����?!������?���(\��?�c��D��?n��w��?�	�Z��?P�$e���?�����?\���(\@��~ǜ?�?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�Ǔ���?�C����?�������?A�ra���?�@۽U��?���Q��?�/�����?�J�LT)�?�������?5�Z(��?XV��?��Q�@�����>�?Po�S3�?!1ogH��?�8Sn�Z�?8Q�H��?�Q���@���
�S�?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?�uS�X�?�P8��?�%m�l��?�I��I��?��������/�X/(�?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?S;>���?�Y���?�gS���?U�j�o�?أp=
��?���tt��? 3`���?���P��?�D�e'~�?�]���?{�G�z@=�A7���?�п�cX�?���؜��?��{�z��?�F��?_fffff�?�F�9���?���S��?��c�0��?k��{<j�?9
�
0�?<
ףp=�?z��w
�?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?r6]����?�������?�	��6f�?���3$��?H�z�G@��S��?XD"���?R��+Q�?$ ����?�#F���?P���Q@]�"�H��?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�6jDRf7�?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?���#�?��t�j�?��qg	��?d���1�?(�)��;�?�������?�O^J��?y�N�?�'��m�?=J�i�?     8�?      @v�u����?"
c���?�[�[�?��
y3�?q�M����?���Q��?�����?evoƃ��?�q�u�?�)���R�?t������?0\���(�?I��p��?q�CZ�y�?)%\����??��"u��?�hJ���?433333����z��?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?[�_�?r���&T�?Vl;!t��?�O��O��?�Q���?0�0q�?�6�)��?7�S\2�?�^�r��?�kD�
��?�G�z�@�o1(��?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?/G�9�?�����T�?`�t����?	�m?���?��Q�@�J��}��?j|��
�?�z�G��?�����?����o.�?�(\��� @�	�x���?+by,Y�?      �?B���?f���?�G�z@�1�2��?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿|�TT�+�?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ�5N�m<�?��2�?�&���?YA�-��?���.�d�?�G�z@O���ii�?%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�<�^�?lq�����?ѭ8��7�?�V8Y+��?��07�Z�?������ܿ]�ڶ�K�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?��;�l�?��{����?��`|��?���!�?@\���(̿Z�S�Ҳ�?�]A6�?��0�:�?A�B)���?7��O	�?�G�z@'�� ��?����?k�_����?��$y���?������?��(\���?��:����?��[y��?�Ў�e��?��^*)�?z^{�?�(\����?�9)�?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���?����/��?~�~��?LgR�L��?|huq���?�p=
ף�?�8G��s�?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?�p��K"�?:�X{��?���.{�?P�l�V��?'��,�?      @���I�8�?�]�L�b�?2&�l�?      �?]|�c���?�z�G�@h��Ơ��?C�Z����?�Nu�w��?��سX��?�R:CW��?H�z�G@�{�͝6�?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�)2��W�?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?��.����?�'#���?�������?&(�iW�?vI�ø_�?G�z�G�?�&A�v�?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?�m�=���?WUUUU��?���a�?v{�e��?���Q��?������?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?l�ģC�?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?��9���?�e���?��G��\�?�����\�?���(\��?:����?Un����?�������?#�R���?]�����?�Q������j;����?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?t��Y��?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?������?9�KO���? ���?R-ŭX�?X�,)D�?\���(\@	`��Np�?P@��}�?��k���?      �?�J���?�������?"t�I�+�?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿぷA�?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��?�'���?�*H^�?�����?Oozӛ��?,\���(�?��x~q��?��2MK�?�`�`�?{���K�?�.�|��?��(\���?�٤�I��?�+����?�#�;��?��oa��?��8���?�Q���ѿH����?� �����?r�q��?܌��! �?���[���?��Q��ۿ�#Bt�?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?I��~j��?fo/���?/����?'N`�4��?��3���?�������:T�+���?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?��O�V�?R8�u�?S{���?��,�1�?:�oO�$�? �G�z��S�hz���?��y����?I`�:�?�5G��`�?4h��J�?      п�P�$��?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?�Gq���?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?:r����?@i���?P��O���?�k�9���?��U�^�?(\���(�?�α	6�?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?����?      �?ŵ�a��? )O��?      @�����?�$�vQ�?����?dȇ���?�?2�խ�?*\���(@��W���?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?�
⛏A�?��P���?4 ��<�?(
P�;�?������@�X0����?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�b=��
�?[̽e��?�)`>�]�?i���/��?o��[�?������?G�x���?���#�?��qPt�?���J��?�T�w��?�Q���?J������?����?���a���?Û�P�?�`8wC�?P���Q�?���Z���?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�m�����?W['s�,�?E�JԮD�?��K�y�?��J�[��?r=
ףp@
�#�F�?U[G[��?;�;��?�	v�o�?�a�a�?������@U��A��?h��Ƅ��?UUUUUU�?���t�?     ��?q=
ףp@����k��?�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?O|-Ϯ��?�X�y"��?%'¸Lr�?c�/�]�?,mG8��?�G�z��?�^���?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?T�k���?���1�?��fy��?���N�R�?Wŵ.���?���(\�@n�-���?(1B���?b'vb'v�?s�ӭ��? �R{���?H�z�G@K3$���?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?�Ȳ���?�YĘ��?9��8���?�鑢3�?^��3��?�G�z��?�*ml|��?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?2E�Ĵ�?	��-��?'m�`�?:o1���?hfffff�?��E T�?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?톘��=�?+P�W
��?���gk�?�������?Z���(\�?�Q�rX��?�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=��_��#�?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?կ~_�:�?�SR�&�?}�K`]�?��<d��?w�C�v�?���Q�ο�*UۄP�?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�??4G0�?������?�~H���?U��oW�?��S�r
�?
ףp=
�?���y[�?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?� �����?{ӛ����?��*��I�?"�nd=6�?������@ }a��?e�F-��?�������?���:%�?V���g�?ףp=
�?´�z�)�?Xe�6�?
ףp=
@�3��x�?�D�Z���?(\���(�?2�b���?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�X�!)b�?��h�D��?��P��9�?�1$0��?}��O���?833333�?&~��.w�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?əPB�?��.���?gL0�h�?l��(�?ףp=
�?��m��\�?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?���|�?      �?��`��?iiiiii�?{�G�z@�iյQ�?\�����?�3�u�?�d�yv6�?f����?���(\�ҿ���#�?�Ұ���?      �?�]8���?��6Ls�?=
ףp=@����a�?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?���-��?�������?�p߃���?y����?hfffff�?fd-c��?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?���1�^�?\	# ���?�߈��?Ľ9�X�?и[���?\���(\�?b�����?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@yU�٬�?T�.�n��?�-�׮�?H{����?������?P���Q�?��/>�?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?
��\���?��\AL��?)us�?      �?433333�?@�����?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?����?CBq�n�?�M���?ABЋf��?hfffff@?��n���?5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?����?�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�5�����?�m�02��?;r����?���	���?����<�?��(\���?�ca�M��?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?E��.��?5�\�`��?���nD�?P��n��?�(\���@v5�/���?�徦�<�?�\AL� �?      �?�������?��Q��?�A���?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?�{Q5��?K�^�/�?(✭��?.�, �y�?!z|��?R���Q@�
"^���?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?s��&�?(W�7�?���xW�?B�HV��?��(\���?�LGuk�?��]���?[�[�@�{�q�?.q����?���Q��?�@����?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?9�m�.�?C�oB��?      �??��(b-�?b�1`�?433333@��
�f�?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?�83���?�{Nm{�?�F�� �?�������?P���Q�?1l(�?9��%*�?�J��?N�J2�x�?*08͸�?hfffff�?���=��?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��76�?�{����?�Pd����?�{c����?�������?���(\��?�ֺ��	�?�r*��?z�Ha��?��R����?�{mĺ��?���Q�濧�7�jq�?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�?wJ��L��?S��?�p���?�������?
ףp=
@�9e���??d~-��?�u�����?����2�?� ?7��?      �?��Ld��?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�z����?��e!&�?�ydF��?�Wt����?*g���?      @�Z�����?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?X���A�?������ @<�z^��?C���,�?�������?\��陌�?�h<*�?�؉�؉�?G�YH_�?�˟�Ѐ�?��Q���?��-�7�?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?P�����?UUUUUU�?�k�1���?O�n�	�?��Q�@$��t�?�e�:�	�?Dy�5��?��:cc�?�b�X,�?
ףp=
@�j��s��?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?5�T3�?233333@牫;X]�?�������?333333�?��W7�?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?M\=���?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?(� .b��?�k�S��?��F����?���w���? �G�z�?�&ɢ�X�?��aJ��?��˝��?�D�y�?�$���?���(\� @��p��A�?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp�\��E�%�?�}��?       @j��_�?��¯�D�?�(\����?0-�+�?d�.���?O��N���?�UfP�h�?];0���?q=
ףp�?�⿞��?�r��Φ�?�n�l�N�?0��x��?3m���G�?|�G�z @�du��x�?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?����-�?��L��L@;K�*�O�?��
��?�������?��R{~��?2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�V����?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?���A��?�RkJ �?j��i���?��Ť��?�����?333333	@�e��O��?U@�'��?�x+�R�??dM2_�?�(S�\��?�(\����B��e��?�9ɻ�	�?     �?vc���?�;�Y�?q=
ףp�?�e���C�?%�����?*��RJ)@f|��O�?D0��fa�?�G�z�?����խ�?u��=M	�?�ڧΪu�?f>����?: 2ܫ`�?�p=
ף�?J�)f�?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?*����Z�?w��{���?)�b���?z9��E�?�0��=)�?�������b��i"�?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?�0�����?      @�	h�l��?t�E]t�?�p=
ף�?r��j4a�?u$_U���?7NӫT�?\:CU��?F�;�5�?433333@E����?����?      �?eK'b���?"�!�!��?������@��Ѐ���?�ao�2 �?�Λ�~b�?����?H݊ÿ�?���(\�ҿ3=�Jg��?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�M���?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?�M�2�?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?:��]��?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?R�p,C.�?������?��U�	��?n��x�>�?��Q��@���Ol�?-����?ӟ���?���;<�?�׷0���?�Q����?���e���?�,B�N�?�
��v��?�߾���?������?P���Q�?z��V��?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?L�Q���?����S��? 0 ��?4և����?433333�?�a����?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?����g�?��r���?\��[���?�4�.��?2}~k���?��Q���?���q(�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�Y��.�?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?���p9�?�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿�_�Be�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?u��׿�?�����?IM0��>�?��I��?�h�k��? R���ѿ��B+���?��M1��?�%�8k��?�C���?�������?P���(\�?~Dk���?Z�yv�<�?��a�
��?��ࣹO�?:&߭��?��Q��@ ah���?�5���?@7���$�?h/�����?�������?�y;Cb�?��j�G�?u�5�o��?���d��?�~��?�G�z��?\�o�nl�?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?[�>���?vP�I��?E8S8B�?������?�5��P^�?����������(�?!ml���?�9�n��?Ѕ�	���?��'q��?�p=
�ӿ�}G�?/������?�k��%�?���g���?8S����?�G�z��� ���V��?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?����*�?)#�`��?��@�x�?�gL���?أp=
�@��ϔ��?��=O�?M4�DM�?���2��?�ܛ���?
ףp=
@������?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?x��l��?Ɏ �U�?�˴�`��?��N��?`���Qؿ�zz����?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�vף]��?L�|9��?m���X��?�B�q��?����:.�?833333�?����?�N"H��?����?Hx`2��?��r:���?������@�P	�_�?
��Y0�?�G*;�?      �?������?��Q��?�-�����?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@��Y���?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ��Ҋ��?�C�>'��?q�l�:��?��'pw�?��
[3�?��Q��@�2����?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?9�߽9&�?(��qg	�?��K�y�?d}�OG��?���Q��?��5Pӹ�?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?W��{3H�?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?<�b���?����?�Pp���?Ŕ��%�?�p=
ף�?�����?2�7���?���A�?���i���?_7��T�?R���Q@yJA���?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?�����?�NϦ�k�?�Ė��w�?���BP�?ףp=
@����?/��Q��?��8��8�?�Z�_�?�������?@���Qȿg9gD�?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��A��?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@C���P�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?���+��?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ʞ2����?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?LG�3�K�?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿR��-�?Шx�?jF���?������?�.�?��?�z�G��?��2}��?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?���@9�?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?      �?r+�z���?9�0s�?�~��i�?s�p5��?�G�z�@ݳ +���?O�TE���?�(፦@��x�b�?��RJ)��?�������??3�/D�?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?���V��?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?i�*�H�?*q4|��?J�J2�x�?���u�	�?���Q�@����W�?�c��)�?c��4�?�.fxx�?�Ŗ����?������@�J}A^�?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?W��#�^�?��I��?      �?	)�L��?ڟ�!T�?��G�z����8I;�?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?��~���?�_��!}�?B�j
��?��XK�?      �?B9=�_��?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�����?�qV��?�z�G��?�	ϻ���?J��I���?�G�z @��w��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?lt�&��?:+��?NB�3�?Ci!��?r�q��?Y���(\�?��F�#�?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�\��f��?ŷ)�N�?����{I�?�����?�N.�E��?��9�
�?R�і�f�?}m���?�t��ap�?��Gǥ�?!q��?8����?�i2�Ɍ�?p�E4��?��(�0��?b�uB���?�j)t�?��
~&�?���gS�?,Ƃ�	��?��0�|l�?����Y�?��jl��?A���5�?z����?րaG��?05����?�{����?�yQ�$�?$K�_0�?&���?ZM�����?��s�x�?WU���?$^�?��?����}��?�f=2��?=�+����?2�լ���?������?�FF�)�?�刲�f�?�O�2��?IYr��7�?a�,q�f�?���ӪY�?4)��х�?u��Y�@��C���?�q�d4�?g�����?��b�?�mkd��?�X���@S�E%;�?�G��6�?��)��[�?�T�b�]�?�~�<�s�?C�[��@�,R��?v���C�?6�Ţp��?�j�1�h�?�ъ�Ka�?(P>$@�~�[RJ�?��|���?Y��>�$�?Oi�l�?��OV�?�="��@�h,����?B�+�?�~����?,e%��a�?��K+���?�U��Dg@�Iʠ��?S[����?83�c��@�c��?�,!�y�?���Wۮ�?�t����?gZ�P��?���ɯ @�
}�p��?o�s<��?"{�֣��?o�!��?�X����?G8�~@8_��\�?�UPa`��?�������?��l.9G�?JierM.�?u(�̴�?��p�]��?8�pq���?Ӕ*2R5�?8� �?`fX�)�?a`���5�?@j�C�j�?v q<��?��=М��?+���c�?��ڕ
�?���ea��?�V�3��?Y|άd�?�>��/��?T4r.�	�?9�M|�?�:�ìw�?d��Ы�?�7;��3�?���f�v�?2:�1�P�?����?��Sfr�?�J<��?�\/�3�?q����?5��5X�?ߌc�
�?9h��s��?�WV�?��߈���?��1��?J�zΤ��?�Wh!��?l�)+�?��튰�?&W�՛�?�9�^S�?�4Ff|[�?��i��?�ά챫�?P���-��?#��**��?��'����?Tp��.%�?iH�x���?�A�k��?M��r��?-��fD�?*�|�$B��I��;�?6����?J�ԇx�?D�p���?��&�<��?RW5u��}u��c�?V�F��?���}���?U��NQ��?S����?I�wJ�z˿*U|�;��?�'�d��?I*����?�]+��O�?�ߒ"��?�ۣ���п�7����?1%��� �?���!��?*U��ʼ�?�^�Iv��?5���?u�I���?�P[�9�?d�r�F�?�1�~��?�L�U���?���=,g�?�O�O��?lP
ۃ�?�
�V�]�?���׺��?�p����?0�8���?�!�����?�Q۰���?Lb��"�?9[��
��?��Z���?X#/�����]6�q5��?��"���?����\�?������?/9-}��?���j���I���-'�?�[\����?v{Z38�?���[<�?�ꆏ�\�?ÕT�ſ���c���?�t�A��?���oU��?J}t���?��~t:x�?T��'����lՎ��?�/5���?�f.O��?P���8�?e����?=�����ԡ�Ȳ�?j&v��?�{ƈs�?�ᇳ�n�?�9͡k��?���8l�?b�M�[��?�+�8�*�?w
X�^q�?˥=�yx�?�"��I��?�����R@1������?�%�61�?B�Z@�+�?�U�x�?���|���?M�{�P�@%��S��?HVu]�%�?w���zd�?�����?�x��?O��2	�@M���=�?;UP �E�?i�@�Vz�?�\�x�?}����?����@�Q+�6�?�)q�?�?��DN'c�?�-v��x�?1_�?����@������?���E�?S,����?6ք\x�?��xL�A�?�j��:=@����E��?`�&�|�?s�Wu �?5Kx�hx�?�Y�c��?�6�x�5@<�<�7��?��b�C�?\��	���?:z��?���7�B�?��-�@L ,�I�?�!��r?�?�K�VS�?��2�j\�?���0���?�Ѻ��@�ؚtZ��?x�Y�>�?�p��\�?�`��Y�?�����?������@권��?(�mS?�??�L�_U�?v�1B�[�?������?�`��	@���K��?�t���M�?�N8bC�?��PcΙ�?O�ɨ&�?�)yx)@�nwl��?) �v�:�?M���բ�?
�)xЧ�?O�*am:�?,��E�@N��@��?{1�}�?sIHӥb�?&�zoĴ�?���,���?����+�?[J(���?�S�����?7a	^��?H}�B��?��qo���?4��-Ve�?�����B�?��e�?g��'p�?w��?Zc+��?ǀڈ���?�A�p�r�?��a��?B){���?���.Ӵ�?:(��l��?m��� ��?8��N���?β��O��?xl�g`@�?g֍'Ž�?�m-(�?!ƕ +�?�|.j�?}���s�?gn�eld�?h�o�ִ�?��̇|��?�פE�$�?�42j��?I�O��?������?ɆQ�l��?�Y��w�?oF��4�?o����?T�Vw���?̔gA|G�?��A�XA�?��p�|c�?Ї�Yk�ӿ���#�?Ht����?~�����?T��P��?d��8���?~8��?|տF��(��?哘_2��?�) wZ�?�*,Y��?]�?BD��?dZ���ܿ���sA�?�9k��?�O���?�U��?���2��?���&׿9�	Ɵe�?��'�6�?�b���\�?�LG����?�mp���?���ؿ�	ގ�?_�G�>��?FӋ�&2�?��2"��?qn>(��?I�^g.޿O�?�	�?�B����?̃P���?�`�'�=�?�mo���?n=�֘%�?�a�m��?� ���?�����?]S�}_�?�\T����?���Cd*�?�,���?2M�����?H����?,_�\Rk�?���.��?"��5�?71H����?�E���?�+����?�{��4�? !�<X��?��Ɣc�?�猤��?M~����?��D��?�F�v�?��R�%�?�D~���?H�����?��f<���?[��5��?�D�sUA�??@iS�?�N<���?�
zQ���?r�/���?��p���?��/���?+[��M�?���T�a�?��Z��?�D+&@�?4g��3)�?Ҩ��?���m0�?��2@���?,�K+��?O%�#�?��n���?L�-Ft��?��QJ3�?j�m[�:�?壅�<�?�zM��?���nؓ�?�v#Q��?��vl	��?�l�y�?�� ���?@.�}O��?�Y�y>9�?	���)h�?�{���?d��s�ȿ����D�?|Zi��?T��NM��?N����?�����?�뮬�@~�G����?�Ж59�?;��U��?*��c!�?O���t�?��j�?��]����?�Q)��?+lK���?�d��t��?�9�+��?��i`�*@j�/����?���p/�?a��X	�?�Dj��?�z*t���?J$ ��@���1��?k3���?��D�G��?w�ME��?�5�et��?�t�a~.@�?�����?��G��?I�����?���V���?h|Q�?T�(=w@�����?q{d�V�?���zf�?��\���?�1�T��?�UIlR�?1J`ΐ��?;��Q�?z1_��^�?LŔ;	�?ڗ�t��?����?���m��?�}v�#�?pPp��A�?����?��K>s�?l�����?;$���?Ec��?�U�^N�?&6��B:�?��3}��?c�� �?n�Z��?j�:�(�?�L�� �?؟\~��?R�*�?q�����?���!G�?>�����?Bkp��?���4x�?����l<�?���f_�?��vgxE�?���%~��?�Z���?:�W��J�?fZ�&@��?��Q��@k'�:Q��?
]���?F5N���?�b"���?X�6T�]�?j��k)j@�4u��?N�,
<�?�*⒅�?3������?�G��?+NN,P@ E�� k�?r�H5�?F�z���?f�|]�?Z��I?V�?'L�˒v�?�M%" �?��3-�?��E����?T�q�!r�?�S�~��?�;�'`�?�X\�7��?������?��X�Q�?̓����?�ڜt���?�w�=-��%��}��?	��:���?��OV�?�>L����?а�����?~@��p躿'=h��?N�F+��?a������?0�:̹�?�A��P�??���Xȿ������?�v����?�jl��?,�?��?�-6:ل�?��Q��@&:6$���?�9�3��?-`�p��?"dhR]u�? g�� :�?���ڟ@Y5���?�,r��?I�Knpp�?�{��w�?���(�?�}�h�@����l��?G�F�!��?�G�!��?�>/��w�?���q�?0��f�@	�-+��?�F��? �?�o.�X��?�|�w�?"}��\+�? ���@[&��?v0p����?�xE�'�?����j�?�*d�A�?�μA1�?�p1�RF�?9GV���?�p�
!�?�B�R{�?݆Ng^j�?���m�?2M� ��?�ͥ¶�?��a9�?��/i�?�?��'���?�c�l��?u��Ŵ�?��ې,�?,ʑ���?[[�=���?����s-�?�N5�,�?�� ����?��Q�?zҮ�'�? �.+y�?�P���?�h��6��?U8 ���?pSd"�?�x�L�?.M2��y�?ip`5 ��?������?�������?��}�'�?5�3���?74�Y�x�?��t���?��+I:k @#��A���?,g��)�?���$u�?���	x�?Glz-��?����\�@�].�_�?�~����?ܖM��?�D/�i��?���S�?4��?���?�m� u=�?���?(��?�����?x�o���?�B�s���?I��n�?��;`Y*�?bD�~��?p�%����?O��l�?=t�P�?��cp�¿�-ؼ���?d'N���?���y��?�(�����?��҈���?��&�ba�?�;�f=�?s�Z"��?���v�?~�E��?�H�rB�?=��qп������?U`����?ӧ#H�W�?�,�����?6� ����?�9�s���8��/��?�p8}�?��8*}X�?�O�;o�?�Pϋ��?��|d;#�?a���?1K����?SU3��m�?#r��?3�c���? |eπ��?4t�׆��?�z��?�l����?hb��v�?$�3��?_��מ��?T�ͨ���?-l����?OA
���?�\8_���?+�r�u0�?�k��� �?���^E��?��̰�$�?������?�*e�rO�?�sE���?+�T/� @R�@`�?'^#=��?������?6 <��?<��_�r�?h�'@�XV:��?��nX��?h�J�V��?6&qe�q�?4�l=���?�l�Ө@8*�#���?�,x��?��x�<K�?�ft�k�?�I�d��? JqH�~ @����T�?���(�}�?ۖkڧU�?�<�2�?�#w{��?A�a�
@3gO(>�?�!��	�?��O���?��c�kd�?����:��?�m���4@��x��?K��f%�?Sz��jq�??mBJ�`�?�����?�X)I=� @��O��1�?K�<���?��jT��?��=��W�?Mn�}u��?��j
H� @HAc�qI�?�Nnb���?�
i3C�?.;�)0�?�nu�L��?�53��7�?��� ��?B�A7�?�8�u�F�?N`\{O6�?.��Z[��?������?NqU�S��?��%�H�?��$�o��?���(��?f_��?_���:��?��u�r�?��j6���?f���?�߁u���?�i����?WЁ5(i�?E)y!j�?Q��d���?(�o�<r�?RmLo��?���.���?��5�^�?��6�?����!�?�z$ ��?b>�{�?�g)�[��?���u��?�$��?���MM�?&�\�ޟ�?bi���?���Zd�?�3���?a�y�_�?!����?��]p���?��T���?<��O��?�MYA��?.l��k��?�7>�CP�?�te���?T�-��?���N���?�4����?mPt߀��?Z��d�?�����?O'���?R�p��l�?a��Gr�?�uk��?㳫$N��?�Uq#�]�?�;y�ފ�?D����?*I�
�B�?�n�/{��?�% m��?��L`2e�?����w�?DƇ��?����� @�(x���?�����?�Lh=c��?���hxw�?Y�����?�d���w@p������?:�TP���?EEb�٢�?�T����?iz'r��?�q>�i @�����?Dcl���?*k,��?8�Q�?�]x ���?�}�j��п�ɛ% ��?��#+���?H۹½�?���
D��?ߝ${��?����K˿�d���>�?.�&����?���)`�?CۡAXj�?Ն9����?��^��C=ߘ���?�R2���?�;KEU��?B��J���?&!��w�?�g')h`ʿӦ�q��?#&k��?���Bz��?s��r�2�?}(��"�?QL���ʿ٦@��?J�8¡��?�آ�s��?_�B`�I�?l�
����?Ak\�.eп^8���?��*��?�npQX��?ڕJ`��?���w1�?�6$��?0<4���?�?T���?�io`�o�?jG�4���?␌�o�?�E�}�`�? P����?�8���?�w����?�/ѻ~��?�%Ȅ���?D@�i��?�bp�n�?-;	�q �?J��u��?
���?E�H���?O�%���? �5�Ò�?a]���?$��g�C�?E��8��?�XK��?J�L�?e�{>��?)AJ�1�?�4W���?q9 ���?��P����?�J8zU�?�x�D���?Д��
2�?U�?����?ht�-a�?ļa�GL�?{�޲_@��n���?_�����?d+����?�-���?��]D�?=�9�G@�IX���?�,��.	�?��X���?�7ۤ�?�v� ��?Z��w��@0�����?^J=vB'�?����[!�?y���s�?�@v�z��?̕��f9@��4�D�?�CP �?q@l"O�?e���?�`���b�?,]���D@#�kw���?k���?������?��֣��?��J�kO�?_EI7@�0�4���?�y��?�,�1�?�����?N,Z�?���X�)�?	� 
q��?��ddW$�?���֝�?P��ꔍ�?�e�6I�?��`X���?��O�^$�?�f.r+�?��I}��?^���?Q����?�����?�l���?�ww��+�?������?�`���?x@�3�y�?������?wH�ɒ��?���y=)�?��^T�<�?�d���?���bv�?yUIlg�?�I�|��?^��}��?#���wQ�?#�5$��?�5a�b�?&_�O�h�?����ڷ�?������?�Si�?�?k���-�?������?ݫ��W�?��9��?/_`�?�R(;;�?�o2���?(f�X�? ��3��?R^K��?�O����?���z��?*\K ��?^�,���?�����T�?�/TW��?]����?GN4��?p]2H��?����;w�?L��י�? 8|��?�����?�S�`Ɋ�?u���g��?M�y�e~�?�CF���?.�q>���?ˋk߳��?]#>��{�?����w��?x�&	*��?m�6���?L�t���?�zK�o��?���h�?�z¥���?��z+"��?a1���?
��M�?��	�y�?�/�DC�?��WE�?$xh�K�?4N3�&�?¥Vy���?�L[�$�?� ��?*���m�?t"���>�?C���k�?�����A�?&������?P ��p,�?��i(�?��X���?����6�?>oM���?�,�����?�UjZk�?lҌ�N�?���V��?!r_�V��?Q�S���?���s8�?�z�(�Z�?z�h9d�?�����?=~e��?�~Y}�?(��\�(�?�]�a���?�$���?�צ��S�?4H�d�+�?Uκ�1I�?�U-}*�?�e��k��?�Q6��?�c+���?.�'#�?�]���(�?�T2V�?o�[��u�?2�����?")Yn��?QO�m���?��#!�m�?E��=���?�f
SI�?ȴ���?På�c��?-�k���?潉&%��?ipp� �?#f)J���?�E.���?��V1��?	WO,�?g?�ۄh�?�����?�Y1y��?���ݮ�?�pC�P�?]��S<��?��Ƥ5�?�������?.�U&��?���w��?ۀ�'x�?�'X7��?�Z�aU1�?�k��	�?���2��?b�LHb��?\o �?"�J D�?5rH��?"PSE��?E�+���?F�`�L��?�<&�T�?ݗ��5��?��/̘��?L���!�?D<|&�v�?R�;^P��?��Y���?q�po$�?Q4I���?�؊F�	�?C���V��? g>_���?�S@u�?Ư�;(�?�����y�?C����?H}����?�>�f��?�E<i�A�?߽��k�?Ѐ@]�?M^W��?�ZJ{fb�?��Њ9�?k�f���?���X�?ǗU�vk�?[�yo�?�I�)C��?7AV� z�?���!��?�?]�gI�?��2�i�?�E���
�?QC� �,�?t0?8��?$��&M��?AA`�/�?��>��?}��D�?�Ar�	��?��>�iy�?���t�?x�i_��?�s��i;�?���/$�?����5�?%�cz�y�?��&<�D�?[Ap�?��?�N����?����g�?����e�?P�b[�x�?��|O@'�?�����J�?^�kAY]�?��ls�?'�eS�e�?�;]~�?ُQ��?ʵWh��?#$K�q�?ɘ8{�?�Rx�I��?z���F��?@��pK�?��~c�?��.��'�?������?�
?�Q��?'&�E2?�?�b�O��?b+\�U�пO�8�?T�?���?��NM~)�?�P=�P��?3���w�?&��uӿ�r:�H��?���t�?��*q���?�$�~�?�-��?����͓�?&�cit��?�����?��i�?<<��?�7�o��?Q��[�?xXV�?9��f�?H���'��?{�ک�?�3>
���?�0c}.��?��I�T�?~�J5��?h����.�?���t���?��/|�u�?�<����?:��s���?��׳��?���D]�?FB?���?�jƬ,��?�3.����?�M_��?��/.��?N�3
���?e(���?8�bo��?�p�6cB�?JF�~��?��{�N�?X����p�?z��Q��?4	L���?6J2�6�?�'5Gze�?޸�4���?O^��Z�?t�����?,]2�I��?�k���?c�+`f6�?I���U��?X	�?���?d�`��?��I����?��૦��?-N�0��?��s��?�h2%��?��;@�-�??�����?�o�$��?n�o�?�A$&���?	i�^A-�?(4n��?�p�qi!�?�q�;���?���r�?&�8�"�?�����?/�ɾ���?�w?�&�?أp=
��?�����"�?I�'(��?ǙA����?��n4���?g�}����?YEiP���?��S��?ml���?kw=`"��?���2�?�Z7�X�?�E���?b��^�$�?2�ʙe)�?��	
3�?���fj�?��ѵ��?�?ܷ��?��S;�`�?�����?�dn����?�n5'P�?r
��(�?��C����?�suJ��?1�k,��?)��>� �?8J�UR��?�]N����?أp=
��?)�����?� 7I"��?)�|i��? ���,��?�#���B�?��|���?\�4����?�����?M%MMv��?֩}���?o��r�6�?�$�$�l�?낉����?ҡI�h��?y�S:Q��?�L��O[�?v~O��E�?�c�l@�!�����?���-��?(�{�z�?	Dĥ)�?���w�?�h�k�?i]����?�G�
!��?�.��U�?5�E���?�SI.>�?��U�T�?܀����?~�{�R��?�|m���?v�����?MF�x
E�?�..��V�?�#�$��?^ �X��?�v{�hb�?�������?8�xJ�?���4f��?�7y�i��?�/�V��?
��s-E�?�d����?]B�,�?B��,�?6�nQ��?��2�r6�?����gq�?�����g�?E��f���?I�Bi��?���^wQ�?`5^k@�?I�{����?W\g��b�?\��&���?��T����?qT�d�?�o'ר�?"';���?�D�qF��?��8����?7�����?�8*݊�?_o�X���?�d3�0�?�DJ����?|1���x�?L�M8^��?of4���?�X\Q��?z�cI��?p�K���?������?E��I���?��I�?�8�2��?o)���?i�=���?*~D�N��?K
M���?�b��[`�?pe�k��?pf��2�?�P�!��?�`�<�#�?�f�9�?�Z+!�?Чӆ��?�<�n���?}YP����?e���v��?���n@�n�A�?!?V����?���%���?�߄�-��?Ѵ6Q#��?z]ُn{@Y}��9��?�=5ɋ��?�Ј��?J�|���?�Z���?L�|9�@m�	P��?�e'��&�?��5�?ѡ�`E��?a�m~w8�?y�4��@q�����?�N~�[T�?��#l�?KZ��(t�?���[�?�� �@���U�?������?�%~u15�?>����@�?�"�6N�?:&U�:@��F�o�?~u��1�?D�V�/�?�+& ��?��[��.�?/��@jq��ͺ�?y�k1M�?�����?�qQ�1��?B����?v��tQ�@�'����?���Iީ�?J�M��.@0���[�?l5�e��?H�����?s���*�?Fx���?×]�@@�ps�/��?심���?������?�wIJ�?��r��?��c2C@yW�6b�?�a�W��?�cC�M�?Y8���I�?�k)��?bf��J@�g�#-�?I�'���?�������?�[0&A^�?�uEʐ��?竍�F.�?v���;�?HI��c�?��b9rC�? Z,���?�����?�սˡ��?٥�E�?ڎ����?|0��6�?��(!H��?	�g����?�=����?�	�9F3�?�`w�?�T����?������?!�Ym�?3���uD�?1���{�?j�Hǣ�? )\����?��#���?��T���?�_ǃ]��?e����?:F0A���?W��X��?��F�Z��?���� �?��f(��?:�l�U�?_Z�9�?��Q�(��?.R)�>h�?P�ɅU�?w]7w,�?�t](��?0�k�h�?�a�����?i���N��?��N��*�?��ڹH��? 4S��?KV_�X�?&^�*3�?�Z�<�q�?w�*��?0;�N���?>C]���?fZ�v�?�{-	�?���.se�?J���?aa��6�?�q�8Ƶ�?{���<�?�Kj���?�BuNJ�?f����?⩩Wz��?H}Z���?�q5h.�?[5f����?G؏�|.�?�;1!�?�0�"oI�?8�թ�?m�$���?�Ϩ���?��O%���?5�&8a��?lz��>��?H��c��?��M�>�?�?C[�� @
lЇ ��?������?�Pb�v�?!˖E�.�?��e���?�UjP�}�?�YV.���?a�]�	�?Y�PMg��?�Fҭ���?�س{X��?:m� ���?�Sf^u�?9Me�U��?)��rЙ�?πj��?Hִy���?Ұ<O� @��fI���?H+Pц/�?�bP6���?�A�H�K�?��
'�?��+9�� @|+m\S�?PB9!���?��P�?������?<4� 9�?1KW���?W+g���?+'��B�?�>V�H�?���pd�?᭺�2�?�+��@�ڷ7�W�?;����E�?ժX�?̠�\�x�?����?U���<�@��^�?��Ǧ�C�?UZ]���?�i���h�?��}�b�?_ad��@Lp�#J�?��h�;�?e�CA�?n��=�x�?P>@�r��?��]��@>�e�<�?��+5�?��B�:�?C&�z�x�?y�G�f�?+*�|t@������?����5�?��X��W�?U�C^�^�?�7_�m�?xl��@V.����?�sʤC�?�"ە2�?���x�?6=Jex��?����@q�D}t$�?@ԕܹ!�?+�9���?�6�'���?q��'�A�?.x	gŘ@�n��l�?܆	�p��?@F�׉U�?>���z��?i���?l!�`�@�?"�5�?F�ug��?4xϨ{p�?����w�?j�e#�?���6�@���E��? ZY�
�?�����?N%�T�y�?�}h鳜�?�KH�4�?n5��3�?'ؔkK��?��n b��?��g*�5�?g�@�?�#(�x��?�7\QѾ�?�g�|�?)�Q�Ҹ�?��NGa��?��ƺ5�?��@SZ��?���(7�?o�"ܞ��?�����?���$�P�?�Tcz@��?������?*���9��?��D6�?-�ޚ���?�7��'q�?�07�:.�?RB^	�?��r1*w�?s�RYc$�?m*����?P0�bs�?��ה�v�?�P b��?�L����?/�����??>g�Z1�?�JУ�?
������?�N����?�]��$�?����3
�?�<�{�;�?)tꊮ�?���h�@�?�ɲ]�&�?/ m 0��?�<@)�
�?������?=A�8���?7(ej>�?]�t���?O·��?W,�����?|�[)�?��/����?�-B�|H�?_#�f��?�'d_��?r��7��?�i�Q�?�Ԉ���?�Sc4mE�?���O]����2m�?V�-��?:��lM�?�d�Aa�?o���?�N��~���i��][�?�5�����? $)h��?hA ���?�Go�'6�?�G�W�� ��2�?b�����?9u#J	�?+hv�
(�?uE�1��?�T'
eH�?�.Bg��?�m����?�d�d��?$��Ԃ�?���a_�?[�f��?8�/v�?��P$	�?١����?:W�z�?��ڸ��?+��\`�?��X#o1�?�N88���?���W,P�?	����y�?�T�(Ŗ�?�;{x���?Ԏ�hi]�?�z)�?�R����?�S�T�y�?�Kx���?�� }���?2��84�?�i�����?[�cǨ�?���/�{�?��%�~>�?���XV�?F3�)Z�?��u����?
���o�?��.��?(S����?�8�&mC�?w�
�m��?��S�$�?ܪX�{�?��_Ș��?���Np�?v��Z��?��k*�?8�?��M7���? �����?~�%��D�?*XʧO�?������?�slg��?�Ҳ^o�?Oq�?��?]�����?�cǇ�z�?1e[����?���=��?#5h���?��V��?�J�2zk�?��|��?����?8��l=�?ND�����?{�k֋�?eJ�2�?�.eb��?_�e��}�?7A��"�?�YEߖ�?K�)G���?��e�m�?;s3�~��?~�qR�6�?����?�4%d1�? z�K��?��g����?��m�?Ʀ�u0��?nV8��?t��T�?���G0��?Ѩj�h�?_v;Z�2�?Hq#��:�?�`��Q%�?J���?_����a�?���&��?��:��?�2��Ѭ�?m�3�?�i�dҝ�?����[��?/�C4��?I�1]h�?oߤ��U�?9s��p#�?a�e�+��?�-_�U�?�+WN���?�"{���?F	�{��?�r�/�?8���$��?��j�M��?{"���W�?X�+�?���.�?����?�&i���?N��?.!o���?�Ix��~�?�&KV��?��:��?�����?Z��px�?0�@���?���
@�h�\��?�ʧ���?f����-�?���#Ã�?6��"�?�7���?���e�?I����?�����?�6;<���?�t�����?/@
��N @�e�)��?|,��z��?�Z퇞��?�K�ц�?T��_7��?+y?ݨ��?`���?`n�̄��?�Y�N	�?a3�Sʆ�?�I��7��?'
���G @�<��	�?�
�aW�?�挛P�?I��[h�?��yGou�?��*I2�?!["7��?����?��W=}D�?�I�P��?;f	C��?�"��E�?@��sL��?A4��?�	�1^��?������?���8��?L��,�?�z�K���?kg�p���?�,���?w1����?�&�OM�?x%�M7�?Q�?�el�?��;G��?�i�(��?MW����?�'�$���?����ְ�?\�Y@�)�?)I���?����ca�?��a d��?�K�Yq��?��Ԟ��?����?��$����?Y�',��?*|�uZ��?�>�pf�?�i%˭T�?��Ymq�?4�����?�0��?S��i+��?�	�;q~�?��@|[��?��B4��?s��G���?2 �|��?������?�ŉ��b�?�S�_Mx�?��/S%Z�?Ba��
�?n�!x�?���|@��?�7�&��?R�1��W�?(����?8�����?��wq!�?���z �?hHE{���?~�B���?�ܺnUV�?0�&G�?+*QK��?�߅[��?�ВW��?��VR��?�P�x��?R9*pT��?�b���?�X4�i�?�֖�?7W�%�?�>~�^[�?�	��?�$����?���?���?n�&��?��,8�?!
d���?Cxdh�?��1�7��?ZEp���?���a_�?�&���?�;�����?W��S�?������?d�&D[��?O�(�Rh�?��?d��?q���X^�?�y�?��x��?������?��Vyԃ�?$GB���?��C?J��?W�~89�?�*5��+�?�}����?Q�3T���?3]U�/��?�CP����?h_�q��?��E���?B�l*n�?�b�kN7�?o��9˦�?tEOqkb�?qEtqFbX
   _n_supportqGhhK �qHh�qIRqJ(KK�qKh<�C}  �  qLtqMbX
   dual_coef_qNhhK �qOh�qPRqQ(KKM�qRh$�B   UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���rN��/a�UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���1��{�UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���Og�.X-��UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���UTWQ]���Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@n�eyp@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@�����@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@7*D**�v@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@Ⱦ�$ݎ@qStqTbX
   intercept_qUhhK �qVh�qWRqX(KK�qYh$�C�K��~�Y�qZtq[bX   _probAq\hhK �q]h�q^Rq_(KK�q`h$�C^iM��X�qatqbbX   _probBqchhK �qdh�qeRqf(KK�qgh$�C8MN�2¿qhtqibX   fit_status_qjK X
   shape_fit_qkMK�qlX   _intercept_qmhhK �qnh�qoRqp(KK�qqh$�C�K��~�Y@qrtqsbX   _dual_coef_qthhK �quh�qvRqw(KKM�qxh$�B   UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@rN��/a@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@1��{@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@Og�.X-�@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@UTWQ]��@Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�n�eyp�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�������Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�7*D**�v�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�Ⱦ�$ݎ�qytqzbX   _sklearn_versionq{X   0.23.1q|ub.