�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?�z�G�{X   coef0q	G        X   tolq
G?PbM���X   CqKdX   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�C�r�*'��?t�@�@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?�z�G�{X   support_q3hhK �q4h�q5Rq6(KM�q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B@              	   
                      "   '   (   +   ,   -   /   7   8   :   ;   A   B   C   F   H   I   J   L   R   S   X   Y   Z   [   ]   `   c   h   i   k   o   r   s   v   w   x   z   |   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �         	                      !  "  #  $  &  (  *  +  -  .  /  3  :  C  D  E  H  K  L  N  O  R  S  V  Y  [  \  `  e  g  i  j  l  n  p  q  r  u  x  |  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                  )   9   =   O   Q   ^   b   e   l   t   �   �   �   �   �   �   �       ,  B  F  I  ^  a  o  v  y  �  �  �  �  �  �  �  �  �  �    q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KMK�qBh"�B�*  �-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?:M�]��?HA@s}�?g0�d��?��7���?\���(\@Un����?�������?#�R���?]�����?�Q�����ƪ+�K�?~r!�f�?�`(vo��?l��';�?�������?��ԩ/��?AR˔���?JL �F�?�>,��?�������?I��q��?�'iq��?�&��?#�����?�Q����?~�aE�?"�z\��?�R����?I��/�?.\���(�?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?L�Q���?����S��? 0 ��?4և����?433333�?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�G��R�?�`�`�?,T����?�Cv����?���Q��?f�s
���?Y�%�X�?��\��?n�ٰ��? )\����?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?�z3��?������?{�̝{�?I�����? ףp=
�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?�u����?�wK�?��?�ef���?tT����?�z�G��?����?���a���?Û�P�?�`8wC�?P���Q�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿ�0�����?      @�	h�l��?t�E]t�?�p=
ף�?(� .b��?�k�S��?��F����?���w���? �G�z�?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?=������?��f���?O���7h�?���t��?���(\��?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp��T����?Z7�"�u@m�����?����T�?�������?�G����?h�[�t�?`o�3���?C�l����?
ףp=
@�t&����?��(��(�?�^mSz��?g�Bg�B�?������@�G,���?�	����?���R{�?��?�c��?���Q��?��r���?\��[���?�4�.��?2}~k���?��Q���?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�X��S��?      �?Ѹ�U�?1�0��?���Q����g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�D̥�
�?�Zk����?��iz�?���\��?��Q���?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?ϙΔ�?a#@i��?M��d�?��,��?      �?Шx�?jF���?������?�.�?��?�z�G��?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?f��;��?~|`d���?|v���?�������?��G�z�?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տəPB�?��.���?gL0�h�?l��(�?ףp=
�?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?��ix�?M��
���?��3�x�?���c�?x�G�z�?�
�����?���!y�?��S��?�����?������ܿ�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?������?�~H���?U��oW�?��S�r
�?
ףp=
�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��,���?�z�G��?����U��?a���{�?      �?�,B�N�?�
��v��?�߾���?������?P���Q�?�X$����?L�:,��?&����?G�N��?\���(�?5�T3�?233333@牫;X]�?�������?333333�?F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿ,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?fo/���?/����?'N`�4��?��3���?��������T��?��gjƻ�?����V�?�����?\���(�?f��UJ��?�!XG��?�����?����vW�?8
ףp=�:N�1��?G�:y�?Y<�&!�?F����?��(\���?���e��?I��/�?i�(�U�?�VC��?T���Q�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?�qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?vP�I��?E8S8B�?������?�5��P^�?�������"&�H
�?�?�4��yO�?��)��?
ףp=
�?����g��?�]����?P�øW�?v�=H]��?��Q���?����?k�_����?��$y���?������?��(\���?�b�)U	�?�s���?�M�isT�?N1�^�?q=
ףp�?L�|9��?m���X��?�B�q��?����:.�?833333�?9gήc��?�Z$�R��?������?�/��/��?033333�4����?�%����?�J:��?v{�e��?���(\��?F��W~�?��f=Q��?�����?DDDDDD�?P���Q�?�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff���>����?      �?0`z��Q�?'u_�?�p=
ף�?���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�? ��2�?S�n0�?���&�_�?I%�e��?�������?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�? �5�0��?�����?B �Gey�?r�q��?��Q���?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?������?������?�X^o�?��<t/�?H�z�G�?����/��?~�~��?LgR�L��?|huq���?�p=
ף�?�0�1���?��8��8�?S�K�?�s����?@
ףp=�??d~-��?�u�����?����2�?� ?7��?      �?���X �?�\�\�?6#�|a�?>6:8���?P���Q�?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�ۇA�?��*�3��?���R�]�?AA�?��(\���?s����`�?�0�0�?��e�s��?���]�(�?�������?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@����?��R�y�?�����?�s@ڦ�?�p=
ף�?��+���?G]t�E�?X?A�x�?Ӱ�,O"�?�z�G�@."t��D�?]t�E�?N����Q�?�^�^�?|�G�z�?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?^���O�?o��o��@�H<�'�?�X�%��?�������?�S�����?8�P\�?��;^�?M�*g��?\���(\�?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?"K�_y�?���,d�?���<�?jhɬ�?�Q���?��Sr��?U����?<����?w�{��?<
ףp=�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?��zZ �?&jW�v%�?t���?X`��?!��Q��?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�п�cX�?���؜��?��{�z��?�F��?_fffff�?��h�D��?��P��9�?�1$0��?}��O���?833333�? *+C[}�?�������?wk�����?e�&Jvm�?��(\��տ쟜�ث�?�$I�$I�?Q�d�?J��I���?0\���(�?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?T�.�n��?�-�׮�?H{����?������?P���Q�?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?M؜�ƹ�?x�5?,�?a�}�I<�?��Z%��?��Q��@K̂��?�O�պ�?�X��F�?      �?�p=
ף�?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?0.Ba��?.�袋.@�
�l�?haz�g�?      �?J""}��?����;�?jZ��m�?�0�9��?��Q���?�_����?      @����,��?[�o�W��?���Q��?,"�j�%�?,-----�?'狗�8�?�`�����?133333�?"
c���?�[�[�?��
y3�?q�M����?���Q��?�!ފ�?c����?��J%%�?��(\���?�G�z�?/������?�k��%�?���g���?8S����?�G�z���4��Y��?���^��?	������?6���+��?|�G�z�?���~�?9"�P9�?<O�����?!������?���(\��?�qV��?�z�G��?�	ϻ���?J��I���?�G�z @�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?֊�q��?��Z��Z@�K��?#e�����?���Q��?
��Y0�?�G*;�?      �?������?��Q��?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?8����?�gS��=�?�~��H�?�Vi�_�?�������?auȒ���?�v%jW�@��s5��?`����?�Q����?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?c�2��8�?l�l��?�����?T��S���?�p=
ף�?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�'*���?mB1rq��?�DI��?�!r���?�Q����?��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?��2���?���?��</�b�?�ռY͛�?H�z�G�?�p^��m�?tT����? ����?����x�?���(\�
@U@�'��?�x+�R�??dM2_�?�(S�\��?�(\�����h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?`���`��?���-��?����w�?��-�jL�?��(\��ſXe�6�?
ףp=
@�3��x�?�D�Z���?(\���(�?�d����?���-���?_l�9��?L��N���?P���Q�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?X���A�?������ @<�z^��?C���,�?�������?aZ�/���?�p��[(�?9�����?���
b�?�������?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?톘��=�?+P�W
��?���gk�?�������?Z���(\�?E�X9�x�?-��,�?)=��'�?��0���?�Q����?"*����?�q�q�?�s�̫~�?+1��JL�?�p=
ף�?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��H��?�z�G�?G��ֳ�?
݋н�?R���Q@��B\&�?�n0E>��?���L�?2 K��?�(\����??V�)��?_�_��?      �?��B�
�?�G�z�?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?4s���?�����?/z�V�4�?~"����?H�z�G�?�h�(���?����?�3��=�?g�=���?�������?8P��A��?�\;0��?<b���e�?y{�X�?      �?���. �?i�`���@jڪ���?��}ylE�?�(\����?�'=��?��fě�?��Xf[�?���¯��?�G�z @R8�u�?S{���?��,�1�?:�oO�$�? �G�z���6"��t�?�[���?�r�@t �?





�?q=
ףp�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?��״��?Ѻ���@��O��?����T�?���(\��?-����?ӟ���?���;<�?�׷0���?�Q����?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�h<*�?�؉�؉�?G�YH_�?�˟�Ѐ�?��Q���?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?���q&��?      �?�ƽ7�?%Ԑ�W��?�z�G��?�n��?�3_�g��?����B�?`V�4[s�?`fffff���83���?�{Nm{�?�F�� �?�������?P���Q�?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?�W���?{�n��?	sG�h��?в�9��?��(\���?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?��k�<��?�k��%�?^�4�y�?��xN%�?433333�?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?�L���z�?X�O���?��F�{�?!���c��?�(\����?�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?���%�?������??�0Yp�?��ퟡz�?r=
ףp�?
��\���?��\AL��?)us�?      �?433333�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?@i���?P��O���?�k�9���?��U�^�?(\���(�?u�-BK�?��T��K�?��x���?>���~��?���Q��?:����?�5��P�?v$����?;�;��?أp=
��?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?�徦�<�?�\AL� �?      �?�������?��Q��?evoƃ��?�q�u�?�)���R�?t������?0\���(�?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?	�F@�?�����?c�I���?l��&�l�?!��Q��?��/����?���T4�?h�v�Q�?�����? ףp=
��2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�y]>d�?g;>)7�?�Ǭ�NR�?&H-/|�?=
ףp=
@�{����?�Pd����?�{c����?�������?���(\��?+e��R�?pА����?�_P�
�?���譺�?��(\���l,����?gH���?���2G�?v�A����?�z�G��?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�m�02��?;r����?���	���?����<�?��(\���?O�t�N>�?�����`�?TBP����?J���h�?
ףp=
@�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?s��&�?(W�7�?���xW�?B�HV��?��(\���?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?�p�|���?���)��?^�3���?h�J� :�?�Q����?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?�'���?�*H^�?�����?Oozӛ��?,\���(�?�wF�?��D'�?6������?�_�_�?�������?��~���?�_��!}�?B�j
��?��XK�?      �?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?����-�?��L��L@;K�*�O�?��
��?�������?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?"�FU��?�71}�?v��3���?�N�Q�S�?�Q����?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?gDAl���?<e�U!�?��-��?'u_[�?�Q����?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�? Jx5��?�a�a�?�;x��<�?�������?�Q���@T,���?T:�g *�?"�[��t�?7.Hj��?�������?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿ�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?��M1��?�%�8k��?�C���?�������?P���(\�?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�����?)�����?�s�H�?�u�y��?�G�z�?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�uS�X�?�P8��?�%m�l��?�I��I��?���������4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?����8��?��*H�?>���h�?�؊���?$\���(�?erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?�S�����?���NV��?��=��?^���?��Q�@�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?���h��?���{��?k 2-�?b�V�;��?�G�z��?���6���?�w���?zkfkl��?�k(���?      @P��-��?�NV�#�?8��m���?�;�#�?333333@qCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�   (   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM�qPh"�B�  (ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M��b��7�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�*Q"��,<�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�&��CQ.D�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M���M/6B�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�pP���%�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�H�-$���(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M�(ӄ2M(M��6;��a@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@������u@S?�&�i@������u@������u@$'�d7J@������u@�h��Lq@������u@������u@������u@������u@������u@������u@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�C
�����qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�C�f�y�q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�CDW�nz��qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�C
�����?qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM�qvh"�B�  (ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@�b��7@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@*Q"��,<@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@&��CQ.D@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@��M/6B@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@pP���%@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@H�-$��@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@(ӄ2M(M@�6;��a�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�������u�S?�&�i�������u�������u�$'�d7J�������u��h��Lq�������u�������u�������u�������u�������u�������u�qwtqxbX   _sklearn_versionqyX   0.21.3qzub.