�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?PbM���X   coef0q	G        X   tolq
G?PbM���X   CqKX   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�C!O	� �?qG�w@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?PbM���X   support_q3hhK �q4h�q5Rq6(KM��q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B�               	   
                                                             !   "   #   $   %   &   '   (   )   *   +   ,   -   .   0   1   2   3   4   5   6   7   8   :   ;   <   =   >   ?   @   A   C   D   E   F   G   H   I   L   M   N   O   P   S   T   U   V   X   Y   Z   [   \   ]   ^   _   `   b   c   d   f   g   h   i   j   l   m   n   o   p   q   r   s   u   v   w   x   y   {   |   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �             	  
                                   !  "  #  $  %  &  '  (  )  *  +  ,  .  /  0  2  3  4  6  7  9  :  <  =  ?  @  C  D  E  F  G  H  I  J  K  L  M  N  O  P  Q  R  U  V  W  X  Y  Z  ]  `  b  c  d  g  h  k  l  m  n  p  q  r  s  t  u  v  w  x  {  |    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                 	                        /   9   B   J   K   Q   R   W   e   k   t   z   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                 -  5  ;  B  S  \  ^  _  a  e  i  j  o  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �      q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KM�K�qBh"�BPK  ��Zb��?��+x���?� �Y]��?����?hfffff@������?�N��N��?��U>R
�?	f���?�G�z@����?      �?ŵ�a��? )O��?      @u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?Un����?�������?#�R���?]�����?�Q�����ƪ+�K�?~r!�f�?�`(vo��?l��';�?�������?R�p,C.�?������?��U�	��?n��x�>�?��Q��@�p�|���?���)��?^�3���?h�J� :�?�Q����?�RkJ �?j��i���?��Ť��?�����?333333	@��ԩ/��?AR˔���?JL �F�?�>,��?�������?i�*�H�?*q4|��?J�J2�x�?���u�	�?���Q�@XD"���?R��+Q�?$ ����?�#F���?P���Q@I��q��?�'iq��?�&��?#�����?�Q����?���|�?      �?��`��?iiiiii�?{�G�z@~�aE�?"�z\��?�R����?I��/�?.\���(�?j|��
�?�z�G��?�����?����o.�?�(\��� @G�u���?�t��6�?ZM��W�?�ɵ��?gfffff@��{G�?����S�?Y�_��?�����B�?֣p=
��?���[�?����NB�?b%c�r�?����]�?hfffff@P,��v�?�������?4:�$�x�?�%����?�G�z�?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?9�߽9&�?(��qg	�?��K�y�?d}�OG��?���Q��?T-����?UUUUUU�?L�5���?�������?ffffff @L�Q���?����S��? 0 ��?4և����?433333�?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?_^MiK��?�q�q�?P����?@�wܛ+�?\���(\�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�4��
:�?(6$�)G�?(��J+z�?v��4��?���(\�@a�B��?�������?' Z�u�?�����?���Q�@�]�L�b�?2&�l�?      �?]|�c���?�z�G�@��U�;�?�ϽF�d�?&���g��?�be�F�?)\���(@�G��R�?�`�`�?,T����?�Cv����?���Q��?f�s
���?Y�%�X�?��\��?n�ٰ��? )\����?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?��S3;��?ĸ_�T>�?��a8%��?�,�י��?q=
ףp@)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?�z3��?������?{�̝{�?I�����? ףp=
�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �?!��m#�?r�q��?�_پ%T�?"Y�B�?{�G�z@S\�C{��?5�rO#,�?64�����?�|�G�j�?ףp=
�@�O�C���?y�5���?�V�ޑ_�?%���^B�?=
ףp=@��n9�
�?�Zg_D��?_j�P�?r1Bm��?H�z�G@�����?�MA�1�?I �����?,|L���?�(\��� @}9�ot��?d����.�?֐��<�?OP�?�z�G��?9��%*�?�J��?N�J2�x�?*08͸�?hfffff�?U[G[��?;�;��?�	v�o�?�a�a�?������@�u����?�wK�?��?�ef���?tT����?�z�G��?����?���a���?Û�P�?�`8wC�?P���Q�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿ��X���?l۶m۶�?�r/js�?]t�E]�?���Q� @�wF�?��D'�?6������?�_�_�?�������?EÓ���?�����?�&z��V�?WUUUU��?���(\�@��e!&�?�ydF��?�Wt����?*g���?      @� �9�$�?h���Q��?�3�s�?�B#�E�?��Q�@�0�����?      @�	h�l��?t�E]t�?�p=
ף�?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?u$_U���?7NӫT�?\:CU��?F�;�5�?433333@]��{��?�����?Iy���?E�,V!�?�Q���@=������?��f���?O���7h�?���t��?���(\��?��O�?�\��\��?��_[�?fC�V�?���Q�@�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?�T����?Z7�"�u@m�����?����T�?�������?� �����?{ӛ����?��*��I�?"�nd=6�?������@+by,Y�?      �?B���?f���?�G�z@��~���?�_��!}�?B�j
��?��XK�?      �?���m,�?שǳkF�?�8��y��?@�Z���?�(\���@�t&����?��(��(�?�^mSz��?g�Bg�B�?������@y�-[Y�?�8�?'�8����?%���E�?�G�z�@��B~���?ƶ#e��?-��k4�??&ǒ::�?{�G�z@
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�G,���?�	����?���R{�?��?�c��?���Q��?��r���?\��[���?�4�.��?2}~k���?��Q���?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�X��S��?      �?Ѹ�U�?1�0��?���Q����9vZC��?X7�"�u�?A ��X�?ƃ'��?�G�z�@�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?%���y��?a8B��?�!!?�Z�?���q6�?<
ףp=�?�D̥�
�?�Zk����?��iz�?���\��?��Q���?����-�?��L��L@;K�*�O�?��
��?�������?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?������?�5��P^�?lN�b�Y�?���v�?�G�z�@�_�0�?�������?|/�����?��Jj+��?
ףp=
	@�@����?�����?���Q{�?(������?�p=
ף@ϙΔ�?a#@i��?M��d�?��,��?      �?Шx�?jF���?������?�.�?��?�z�G��?��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�?"�FU��?�71}�?v��3���?�N�Q�S�?�Q����?Ŀ�y/��?.V�oD��?0�Է�N�?]2�h��?ףp=
�@=��a��?}T$;f)�?�|��O�?�UO���?��(\��@f��;��?~|`d���?|v���?�������?��G�z�?�9ɻ�	�?     �?vc���?�;�Y�?q=
ףp�?�����?IM0��>�?��I��?�h�k��? R���ѿݘ��2��?      �?)�gf��?B7%�!6�?��(\��տəPB�?��.���?gL0�h�?l��(�?ףp=
�?�YĘ��?9��8���?�鑢3�?^��3��?�G�z��?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?��ix�?M��
���?��3�x�?���c�?x�G�z�?�
�����?���!y�?��S��?�����?������ܿ��=�9�?�[��"e�?�+U��R�?�Gq�>�?��Q���?\��Z�?�$I�$I�?��ԉ#\�?����>4�?]���(\@�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?������?�~H���?U��oW�?��S�r
�?
ףp=
�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��,���?�z�G��?����U��?a���{�?      �?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?�,B�N�?�
��v��?�߾���?������?P���Q�?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?5�T3�?233333@牫;X]�?�������?333333�?Za�T�
�?�1���N�?D��car�?�MҷV��?H�z�G@�,ۈO�?.�q˸�?4-�����?O�0���?Y���(\	@F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿ,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?�T��?��gjƻ�?����V�?�����?\���(�?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���e��?I��/�?i�(�U�?�VC��?T���Q�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?��<���?      �?��(�r�?��a	G��?���(\�@���<�+�?e�/��b�?>�t�Z�?X,
�?R���Q@{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@��=Qr�?7r#7r#�?y�sJiM�? ��c��?433333�?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?vP�I��?E8S8B�?������?�5��P^�?�������"&�H
�?�?�4��yO�?��)��?
ףp=
�?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?B(w}1�?p�j:�?�ⷆX��?�H1�_��?���(\�@����g��?�]����?P�øW�?v�=H]��?��Q���?����?k�_����?��$y���?������?��(\���?�b�)U	�?�s���?�M�isT�?N1�^�?q=
ףp�?C�oB��?      �??��(b-�?b�1`�?433333@L�|9��?m���X��?�B�q��?����:.�?833333�?�_�^�/�?      �?K��>�?0�9�a�?������@��Lf�@�?�!��uy�?������?�aS���?�G�z@Eb���?��Y@�H�?�|��X.�?�������?��Q��	@�4����?�%����?�J:��?v{�e��?���(\��?�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?�_����?��.��@�ʌ����?�v���?��Q���?���Y�?�	g�	g�?ya��w�?!s��2�?�p=
ף@�>����?      �?0`z��Q�?'u_�?�p=
ף�?i�+s�?333333�?`�>��R�?��.���?q=
ףp@�*�N��?
ףp=
�?_�6�?:����R�?�p=
ף@���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�?��L��?�q�q�?G`3�!�?O���t:�?R���Q@r	����?�8��8�@�m��D�?�O�?���?ףp=
��?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?|A� *��?�袋.�@��k{�?W�+���?H�z�G�? �5�0��?�����?B �Gey�?r�q��?��Q���?yϠ�%�?      �?^���т�?      �?�G�z�@S;>���?�Y���?�gS���?U�j�o�?أp=
��?EtA%�?/���}�?�f�M��?��¯�D�?���Q�@�(ؚ��?�{a��?Vu�o� �?      �?��(\���?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?������?������?�X^o�?��<t/�?H�z�G�?��=O�?M4�DM�?���2��?�ܛ���?
ףp=
@2�7���?���A�?���i���?_7��T�?R���Q@�0�1���?��8��8�?S�K�?�s����?@
ףp=�??d~-��?�u�����?����2�?� ?7��?      �?����?      �?eK'b���?"�!�!��?������@���X �?�\�\�?6#�|a�?>6:8���?P���Q�?%�����?*��RJ)@f|��O�?D0��fa�?�G�z�?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?%n����?      �?7��S�?��/���?�p=
ף@�m�=���?WUUUU��?���a�?v{�e��?���Q��?�@��+W�?��)o���?�߾���?      �?������@�ۇA�?��*�3��?���R�]�?AA�?��(\���?�ӄ���?R���Q@���K���?����*��?�(\����?s����`�?�0�0�?��e�s��?���]�(�?�������?�@�,��?I�$I�$�?x�?q�?u<@�La�?\���(\�?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?����?��R�y�?�����?�s@ڦ�?�p=
ף�?��+���?G]t�E�?X?A�x�?Ӱ�,O"�?�z�G�@�n���?H���x�?6?�x�o�?�#�	<�?R���Q@��;�l�?��{����?��`|��?���!�?@\���(̿�����?�NϦ�k�?�Ė��w�?���BP�?ףp=
@�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?p;̞��?      @�њ�%g�?'u_[�?�������?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?^���O�?o��o��@�H<�'�?�X�%��?�������?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?�S�����?8�P\�?��;^�?M�*g��?\���(\�?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?�}��?       @j��_�?��¯�D�?�(\����?�aݚ
�?(������?� R�M�?��7��M�?       @"K�_y�?���,d�?���<�?jhɬ�?�Q���?�-J���?���|�?�o�vE��?T�P�B��?�G�z@��Sr��?U����?<����?w�{��?<
ףp=�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?��zZ �?&jW�v%�?t���?X`��?!��Q��?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?��[y��?�Ў�e��?��^*)�?z^{�?�(\����?�C�>'��?q�l�:��?��'pw�?��
[3�?��Q��@�
⛏A�?��P���?4 ��<�?(
P�;�?������@�'#���?�������?&(�iW�?vI�ø_�?G�z�G�?t� %��?.�袋.�?����2`�?��H	9�?=
ףp=@���?�m۶m�@��X)�O�?�\.�?)\���(�?�r�4�?�;�;�?ڡf6�K�?�s�9��?�Q����?t}ja>o�?\�-�=�?�Jpv��?��|j��?������� *+C[}�?�������?wk�����?e�&Jvm�?��(\��տ�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?P�����?UUUUUU�?�k�1���?O�n�	�?��Q�@t��!���?,�X��?^*��U��?�:�>c�?��Q��@*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?Q�����?I�$I�$�?���Y�?z��!y�?333333�?����0��?�x��ܷ�?Y1"�	l�?l#֥���?��Q��	@��#���?�rcˍ-�?���'��?8��{�?@�z�G�?/9(��?.�袋.
@�*����?�������?�������?{��*W��?     @�E!��p�?�$I�$��?�G�z��?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?0.Ba��?.�袋.@�
�l�?haz�g�?      �?J""}��?����;�?jZ��m�?�0�9��?��Q���?�e�:�	�?Dy�5��?��:cc�?�b�X,�?
ףp=
@��(��?7�Y�"�?ޤ�=%�?{�!���?���Q� @�_����?      @����,��?[�o�W��?���Q��?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@,"�j�%�?,-----�?'狗�8�?�`�����?133333�?"
c���?�[�[�?��
y3�?q�M����?���Q��?�!ފ�?c����?��J%%�?��(\���?�G�z�?/������?�k��%�?���g���?8S����?�G�z��������?�Qf�,�?z�<���?�%���x�?Z���(\@4��Y��?���^��?	������?6���+��?|�G�z�?������?�ol���?})3=[t�?��{a�?=
ףp=@���~�?9"�P9�?<O�����?!������?���(\��?���`�?��`Q�(�?w
R�VO�?�>���?)\���(@�qV��?�z�G��?�	ϻ���?J��I���?�G�z @�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?֊�q��?��Z��Z@�K��?#e�����?���Q��?����t�?���j?�?��y��X�?sƎ�e�?������@��sr��?��3���?�V��?��~5&�? ףp=
׿
��Y0�?�G*;�?      �?������?��Q��?�%��H��?7��<�?zx� ���?]t�E�?q=
ףp@Ũ���?WUUUUU�?%�[P�~�?�������?�(\���@X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?C�Z����?�Nu�w��?��سX��?�R:CW��?H�z�G@���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?E��.��?5�\�`��?���nD�?P��n��?�(\���@ 3`���?���P��?�D�e'~�?�]���?{�G�z@�j���?�B��X��?�����0�?.ܴE�?��Q�@��TD��?x!�����?�x�;���?���&P��?�p=
ף@����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?8����?�gS��=�?�~��H�?�Vi�_�?�������?auȒ���?�v%jW�@��s5��?`����?�Q����?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿ����?CBq�n�?�M���?ABЋf��?hfffff@�%[b�F�?!t��B�?d&�X�1�?��/���?�������?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?:�SR�?���7���??	-zռ�?��y�?�������e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?c�2��8�?l�l��?�����?T��S���?�p=
ף�?Jt_�h��?߈�N�@(���'<�?ZZZZZZ�?�G�z�?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?K�^�/�?(✭��?.�, �y�?!z|��?R���Q@=B�k��?g�K1_h�?;9�=-�?$�D"��?q=
ףp�?�'*���?mB1rq��?�DI��?�!r���?�Q����?F_L�D��?:��8���?�\�]�G�?l�����?������ @^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?�\7z�?���"��?����}�?7�j�?H�z�G@ �X��?
ףp=
�?�Ѣ�ǃ�?�;⎸#�?      @��2���?���?��</�b�?�ռY͛�?H�z�G�?��2�?�&���?YA�-��?���.�d�?�G�z@'�CU$
�?      �?�t�U�%�?.�#EC�?��Q�@�h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?��p����?      �?��e�N�?�������?R���Q@���S��?��c�0��?k��{<j�?9
�
0�?<
ףp=�?Z�yv�<�?��a�
��?��ࣹO�?:&߭��?��Q��@Xe�6�?
ףp=
@�3��x�?�D�Z���?(\���(�?��i�,�?ףp=
��?���b��?,Fڱ�?��Q�@E� �?      �?��ԉj��?��|�nS�?333333	@X���A�?������ @<�z^��?C���,�?�������?�miV���?�U�;���?P�l�V��?A�Iݗ�?�z�G�@aZ�/���?�p��[(�?9�����?���
b�?�������?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?톘��=�?+P�W
��?���gk�?�������?Z���(\�?48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@���*�_�?۶m۶m�?E������?�n���?�p=
ף@E�X9�x�?-��,�?)=��'�?��0���?�Q����?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?h��Ƅ��?UUUUUU�?���t�?     ��?q=
ףp@"*����?�q�q�?�s�̫~�?+1��JL�?�p=
ף�?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?�Fm�}�?�/Rm���?q�Q>	�?ݫ`���?=
ףp=@n��w��?�	�Z��?P�$e���?�����?\���(\@{^Q�h�?       @��Tf,�?�7�7�?�G�z @��*@�?:��8���?�O�Xs-�?���#B�?��Q���?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?����*�?)#�`��?��@�x�?�gL���?أp=
�@�!K���?)^ ���?u�`6�?���j��?q=
ףp�?,$��?>~&.'�?      �?nt<iE��?������@4s���?�����?/z�V�4�?~"����?H�z�G�?�h�(���?����?�3��=�?g�=���?�������?8P��A��?�\;0��?<b���e�?y{�X�?      �?)�>i�??!AF��?�VYo���?������?��Q��@���. �?i�`���@jڪ���?��}ylE�?�(\����?�'=��?��fě�?��Xf[�?���¯��?�G�z @v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@�6"��t�?�[���?�r�@t �?





�?q=
ףp�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�����X�?t�����?�^Y�?��??��5���?ףp=
�?��0��?R�}�=�?ӗYl�n�?.�袋.�?�Q���@�74J�_�?*6\u��?�$8����?�/t���?      @�h��g��?O ���E�?��mQx��?��vY��?���(\��?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?!ml���?�9�n��?Ѕ�	���?��'q��?�p=
�ӿ��״��?Ѻ���@��O��?����T�?���(\��?-����?ӟ���?���;<�?�׷0���?�Q����?m��C�?      �?2zW�]6�?��L��?���(\�@&�6-��?�����?d6�^3]�?��/�R/�? \���(�?ۆ����?wT��~�?�f!b��?���I���?��Q�@���ʦ�?�6f�@��?�~�ϓ�?FM0��>�?�G�z�@d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?P�H �?:��8���?Ta�z`�?�'�����?�G�z�@�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?_�;I*��?k��FX�?e�5���?J����?R���Q@�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�h<*�?�؉�؉�?G�YH_�?�˟�Ѐ�?��Q���?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?���q&��?      �?�ƽ7�?%Ԑ�W��?�z�G��?�83���?�{Nm{�?�F�� �?�������?P���Q�?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?�W���?{�n��?	sG�h��?в�9��?��(\���?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?W����?��8��8�?      �?Au���?�������?wJ��L��?S��?�p���?�������?
ףp=
@�X�y"��?%'¸Lr�?c�/�]�?,mG8��?�G�z��?��k�<��?�k��%�?^�4�y�?��xN%�?433333�?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?�o�����?��%�̀�?�\"�0�?P[AG:��?�(\����?erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?H��O �?���C��?£^b֑�?���;�L�?�z�G�@��S��?I�$I�$�?�����?���w��?�������?�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?~�W�f��?y@�z��?�{b�?�W�^�z�?�z�G�@�$�vQ�?����?dȇ���?�?2�խ�?*\���(@�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?���%�?������??�0Yp�?��ퟡz�?r=
ףp�? '�Q�^�?ᖚ�?C�7�y�?4H�4H��?���(\�@
��\���?��\AL��?)us�?      �?433333�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?����?�N̓���?�[����?*) �'�?\���(\	@@i���?P��O���?�k�9���?��U�^�?(\���(�?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?u�-BK�?��T��K�?��x���?>���~��?���Q��?:����?�5��P�?v$����?;�;��?أp=
��?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?�徦�<�?�\AL� �?      �?�������?��Q��?r�2�F�?�zۜ��?z!I�,�?c[:��c�?�p=
ף@evoƃ��?�q�u�?�)���R�?t������?0\���(�?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?Se�;f�?h����@A�j�}��?�WJ�B��?S���Q @	�F@�?�����?c�I���?l��&�l�?!��Q��?{���T�?=]�΁A�?�DJ#��?���e�?|�G�z@��/����?���T4�?h�v�Q�?�����? ףp=
���_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?����S�?�N�u.�?�&$a��?���7�?      @&1��T��?2w��!�?��WK��?t���1�?433333@2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�=�,;��?!G%޸��?������?ُ�؏��?�G�z�@�Q���?6��<�?@(��?�;�;�?أp=
�@�{����?�Pd����?�{c����?�������?���(\��?�J�LT)�?�������?5�Z(��?XV��?��Q�@r6]����?�������?�	��6f�?���3$��?H�z�G@Sª����?      �?�	*�/�?W�<�?R���Q@&�-ʰ�?�.]�6�?���}���?K��0a]�?������@�C����?�������?A�ra���?�@۽U��?���Q��?L��,�(�?}�>C��?�t��l��?('����?)\���(@l,����?gH���?���2G�?v�A����?�z�G��?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�m�02��?;r����?���	���?����<�?��(\���?���]�?��g����?1sJJ��?��f$/��?���Q�@�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?s��&�?(W�7�?���xW�?B�HV��?��(\���?�|��	�?b�־a�?pA�D�?���rȔ�?H�z�G@�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?����Z�?+�O��d�?���s�?���rD��?������@PPvI�?]�����?ea����?m۶m۶�?
ףp=
@q�ک��?      @���<X�?��=���?333333�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?��]���?[�[�@�{�q�?.q����?���Q��?y��RE�?n,�Ra�?�$\Z�?��S�p�?�������?:M�]��?HA@s}�?g0�d��?��7���?\���(\@¶�F�s�?0w�fs�?)���k�?y�!���?{�G�z@Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?�'���?�*H^�?�����?Oozӛ��?,\���(�?(� .b��?�k�S��?��F����?���w���? �G�z�?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp�^e�NF��?�}�K�`�?GT��a�?&Դ���?P���(\�?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?�G����?h�[�t�?`o�3���?C�l����?
ףp=
@h�����?��1����?�IF��?�_{�e��?��G�zĿ׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?gDAl���?<e�U!�?��-��?'u_[�?�Q����?�X$����?L�:,��?&����?G�N��?\���(�?fo/���?/����?'N`�4��?��3���?�������f��UJ��?�!XG��?�����?����vW�?8
ףp=��qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?��Q����?�~��?O10%	s�?�M����?�G�z�׿9gήc��?�Z$�R��?������?�/��/��?033333�F��W~�?��f=Q��?�����?DDDDDD�?P���Q�? ��2�?S�n0�?���&�_�?I%�e��?�������?�r*��?z�Ha��?��R����?�{mĺ��?���Q�濇���/��?~�~��?LgR�L��?|huq���?�p=
ף�?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�ݭ����?yþ�\�?�CM`��?�w��K�?�p=
��?."t��D�?]t�E�?N����Q�?�^�^�?|�G�z�?�":>ɗ�?���ע�?���'-�?�R71�?      迃ao�2 �?�Λ�~b�?����?H݊ÿ�?���(\�ҿ Jx5��?�a�a�?�;x��<�?�������?�Q���@�п�cX�?���؜��?��{�z��?�F��?_fffff�?G���;�?�x+�R�?gj��?�r4.G��?��Q�@��h�D��?��P��9�?�1$0��?}��O���?833333�?쟜�ث�?�$I�$I�?Q�d�?J��I���?0\���(�?T�.�n��?�-�׮�?H{����?������?P���Q�?������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z���.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?�SR�&�?}�K`]�?��<d��?w�C�v�?���Q�ο(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿ����Z�?r��Z�@� ��r�?g��|�Q�?033333�Ni�3�?�l�����?��+���?�S�n�?!��Q��?��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?U@�'��?�x+�R�??dM2_�?�(S�\��?�(\���࿁�M1��?�%�8k��?�C���?�������?P���(\�?� �����?r�q��?܌��! �?���[���?��Q��ۿ�t�!O�?��+��+�?��\�2�?�2����?`���(\�?`���`��?���-��?����w�?��-�jL�?��(\��ſ�d����?���-���?_l�9��?L��N���?P���Q�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?�����?)�����?�s�H�?�u�y��?�G�z�?��B\&�?�n0E>��?���L�?2 K��?�(\����??V�)��?_�_��?      �?��B�
�?�G�z�?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?R8�u�?S{���?��,�1�?:�oO�$�? �G�z���i����?T����|�?�;x�]z�?,d!Y��?P���Q�?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�?lq�����?ѭ8��7�?�V8Y+��?��07�Z�?������ܿKY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(쿖���8��?��*H�?>���h�?�؊���?$\���(�?�L���z�?X�O���?��F�{�?!���c��?�(\����?�S�����?���NV��?��=��?^���?��Q�@����?��Pp%��?kub�Q�?̟�Ѐ%�?�������I)i���?�{0�I��?KU���?�X�����?@
ףp=⿃�*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?_������?���h��?�����?\t�E]�?�������?���fR�?:�:��?�Pk����?ק�����?��Q�	@���h��?���{��?k 2-�?b�V�;��?�G�z��?���6���?�w���?zkfkl��?�k(���?      @+e��R�?pА����?�_P�
�?���譺�?��(\���u��=M	�?�ڧΪu�?f>����?: 2ܫ`�?�p=
ף�?P��-��?�NV�#�?8��m���?�;�#�?333333@qCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�  O   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM��qPh"�B  !O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� ��� 3#Yÿ!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �!O	� �qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@tF*44q�?qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qG�w@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�Czug	���qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�C��^8��q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�C�<t|�E��qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�Czug	��?qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM��qvh"�B  !O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?�� 3#Y�?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?!O	� �?qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�tF*44q��qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qG�w�qwtqxbX   _sklearn_versionqyX   0.21.3qzub.