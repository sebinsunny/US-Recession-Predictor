�csklearn.svm._classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX
   break_tiesq�X   kernelqX   rbfqX   degreeqKX   gammaq	G?PbM���X   coef0q
G        X   tolqG?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   n_features_in_qKX   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�q cnumpy
dtype
q!X   f8q"K K�q#Rq$(KX   <q%NNNJ����J����K tq&b�C����?�U�^��?q'tq(bX   classes_q)hhK �q*h�q+Rq,(KK�q-h!X   i8q.K K�q/Rq0(Kh%NNNJ����J����K tq1b�C               q2tq3bX   _gammaq4G?PbM���X   support_q5hhK �q6h�q7Rq8(KM��q9h!X   i4q:K K�q;Rq<(Kh%NNNJ����J����K tq=b�B�                             "   &   (   .   0   3   5   8   ;   ?   @   A   D   F   J   L   O   R   S   X   [   _   a   c   d   f   j   l   n   s   u   v   z   ~   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                                     !  $  %  '  )  *  +  -  .  5  6  9  <  >  ?  B  D  K  L  P  Q  S  T  U  V  X  Z  [  ^  _  a  c  d  e  g  h  i  j  p  s  t  v  x  z  }  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                             '  *  .  0  :  =  @  B  C  E  G  H  J  K  M  N  O  Q  S  U  W  Z      *   /   Q   V   \   o   p   |   �   �   �   �   �   �     J  k  {    �  �  �  �  �  �  �  �  �  �  �  �  �       -  [  \  ]  ^  _  `  a  q  t  x  y  z  {  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                    "  #  $  *  +  ,  -  7  9  :  C  G  H  I  M  O  Q  S  T  U  V  W  X  Y  Z  [  `  a  d  g  i  m  n  o  p  r  s  t  u  x  y  z  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  q>tq?bX   support_vectors_q@hhK �qAh�qBRqC(KM�K�qDh$�B�]  :�SR�?���7���??	-zռ�?��y�?�������V�o@��?u�-BK�?��T��K�?��x���?>���~��?���Q��?f[t��?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?���[�?����NB�?b%c�r�?����]�?hfffff@Wd���'�?Qn�p&�?�؉�؉�?�*����?��M�`�?�p=
ף@9�>����?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�?�aݚ
�?(������?� R�M�?��7��M�?       @St��i��?�b�)U	�?�s���?�M�isT�?N1�^�?q=
ףp�?D����?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?0�|L��?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?��j�G�?u�5�o��?���d��?�~��?�G�z��?\�o�nl�?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?[�>���?����=��?|�Zj�M�?������?���;��?�p=
ף�?��"�$��?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?8K����?PPvI�?]�����?ea����?m۶m۶�?
ףp=
@���UY:�?���\�?�^o�?�?Q�/��?^̧^̧�?�(\����?�XrYǾ�?vP�I��?E8S8B�?������?�5��P^�?����������(�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�9��-c�?!ml���?�9�n��?Ѕ�	���?��'q��?�p=
�ӿ�}G�?V�gb�?��W�l��?U�����?_�HI��?�������?��h~3�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?�!ފ�?c����?��J%%�?��(\���?�G�z�?�~���?f�s
���?Y�%�X�?��\��?n�ٰ��? )\����?�b �*�?/������?�k��%�?���g���?8S����?�G�z��� ���V��?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?9�IA�?{���T�?=]�΁A�?�DJ#��?���e�?|�G�z@��F �?�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?��m����?ӏK�K�?��{���?���S��?{���g�?P���Q�?�Z(O,k�? �X��?
ףp=
�?�Ѣ�ǃ�?�;⎸#�?      @3����?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@c-�Gb�?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?P�ϸ=�?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?עWG�?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?K]E!�6�?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?y���t��?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?%����?erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?�J/��?:����?�5��P�?v$����?;�;��?أp=
��?�[9�.�?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?���@���?��a��z�?�����?�5�3z�?H�z�G@������?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@j��!��?x��l��?Ɏ �U�?�˴�`��?��N��?`���Qؿ�zz����?8����?�gS��=�?�~��H�?�Vi�_�?�������?�11�G��?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�vף]��?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?ѳ!s��?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?�h�(���?����?�3��=�?g�=���?�������?���w ��?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?�D̥�
�?�Zk����?��iz�?���\��?��Q���?��е:�?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?l,����?gH���?���2G�?v�A����?�z�G��?fÿ���?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��K�?�
�����?���!y�?��S��?�����?������ܿ����c��?�#tT��?®b�?	�e^��?�m۶m�? ףp=
�?�)�9�?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�<��2��?�N"H��?����?Hx`2��?��r:���?������@�P	�_�?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?It���?"K�_y�?���,d�?���<�?jhɬ�?�Q���?D�&Dq�?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?�-{X�?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?�u����?�wK�?��?�ef���?tT����?�z�G��?��-��?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?s����`�?�0�0�?��e�s��?���]�(�?�������?ApMrx(�?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?'���/��?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?ű�r��?
��Y0�?�G*;�?      �?������?��Q��?�-�����?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?����em�?׊��+��?Y�����?"$�A���?�(\���@K������?F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿr���;�?�&�j��?7��P^C�?F�����?q=
ףp�?��G�z�?:�5+�?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?�~�A
�?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ��Ҋ��?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?�X��e�?���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�?�k�6��?�Fm�}�?�/Rm���?q�Q>	�?ݫ`���?=
ףp=@�+H���?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�Ǔ���?S\�C{��?5�rO#,�?64�����?�|�G�j�?ףp=
�@ �K.R�?9�߽9&�?(��qg	�?��K�y�?d}�OG��?���Q��?��5Pӹ�?�מ���?�i�i�?Q�XW��?�R�~���?      �?t��3��?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?W��{3H�?�y�]��?]�)~I��?��@��[�?�{����?���(\�@#i��K�?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?Eb���?��Y@�H�?�|��X.�?�������?��Q��	@�ڱ���?��t�j�?��qg	��?d���1�?(�)��;�?�������?�O^J��?evoƃ��?�q�u�?�)���R�?t������?0\���(�?I��p��?q�CZ�y�?)%\����??��"u��?�hJ���?433333����z��?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?2�7���?���A�?���i���?_7��T�?R���Q@yJA���?/G�9�?�����T�?`�t����?	�m?���?��Q�@�J��}��?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿|�TT�+�?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ�5N�m<�?���+*�?�-шs��?���ҋ�?�#o��?q=
ףp@N�Π21�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?��;�l�?��{����?��`|��?���!�?@\���(̿Z�S�Ҳ�?/��Q��?��8��8�?�Z�_�?�������?@���Qȿg9gD�?����?k�_����?��$y���?������?��(\���?��:����?��+���?G]t�E�?X?A�x�?Ӱ�,O"�?�z�G�@����� �?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?�p��K"�?뚖f�?1ܫ`���?��Z(~�?�;�;�?@\���(̿O�e���?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?��.����?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��A��?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?��*@�?:��8���?�O�Xs-�?���#B�?��Q���?��;���?�m�=���?WUUUU��?���a�?v{�e��?���Q��?������?�=�,;��?!G%޸��?������?ُ�؏��?�G�z�@������?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@C���P�?Un����?�������?#�R���?]�����?�Q������j;����?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?t��Y��?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ʞ2����?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?������?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?��9k��?P@��}�?��k���?      �?�J���?�������?"t�I�+�?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿぷA�?"&�H
�?�?�4��yO�?��)��?
ףp=
�?�=4Q�S�?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?I��~j��?�����?�Qf�,�?z�<���?�%���x�?Z���(\@��w]�f�?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?��O�V�?�}�!���?��Sڃ�?xE.�;	�?��}A�?��Q�@�=k,�y�?��y����?I`�:�?�5G��`�?4h��J�?      п�P�$��?@i���?P��O���?�k�9���?��U�^�?(\���(�?�α	6�?�$�vQ�?����?dȇ���?�?2�խ�?*\���(@��W���?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?LG�3�K�?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?���#�?��qPt�?���J��?�T�w��?�Q���?J������?����?���a���?Û�P�?�`8wC�?P���Q�?���Z���?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿR��-�?�X�y"��?%'¸Lr�?c�/�]�?,mG8��?�G�z��?�^���?��H��?�z�G�?G��ֳ�?
݋н�?R���Q@X�C���?Шx�?jF���?������?�.�?��?�z�G��?��2}��?���1�?��fy��?���N�R�?Wŵ.���?���(\�@n�-���?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?�Ȳ���?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?���@9�?2E�Ĵ�?	��-��?'m�`�?:o1���?hfffff�?��E T�?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?t}ja>o�?\�-�=�?�Jpv��?��|j��?�������~���-�?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?կ~_�:�?c�2��8�?l�l��?�����?T��S���?�p=
ף�? ���P��?}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@�y��L(�?v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@�����?������?�~H���?U��oW�?��S�r
�?
ףp=
�?���y[�?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?� �����?{ӛ����?��*��I�?"�nd=6�?������@ }a��?e�F-��?�������?���:%�?V���g�?ףp=
�?´�z�)�?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?��zZ �?&jW�v%�?t���?X`��?!��Q��?���f �?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?əPB�?��.���?gL0�h�?l��(�?ףp=
�?��m��\�?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?      �?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?���-��?�������?�p߃���?y����?hfffff�?fd-c��?��mW(��?333333�?"�*|��?���?333333@��K���?\	# ���?�߈��?Ľ9�X�?и[���?\���(\�?b�����?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?
��\���?��\AL��?)us�?      �?433333�?@�����?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�5�����?�m�02��?;r����?���	���?����<�?��(\���?�ca�M��?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?�徦�<�?�\AL� �?      �?�������?��Q��?�A���?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?�*�N��?
ףp=
�?_�6�?:����R�?�p=
ף@}�"�>�?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?s��&�?(W�7�?���xW�?B�HV��?��(\���?�LGuk�?��O�?�\��\��?��_[�?fC�V�?���Q�@��8܅�?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?�_{��\�?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?�83���?�{Nm{�?�F�� �?�������?P���Q�?1l(�?�$�@�?      �?i|�NT�?칊e��?�G�z�?�����v�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?���V��?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��??d~-��?�u�����?����2�?� ?7��?      �?��Ld��?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?�h<*�?�؉�؉�?G�YH_�?�˟�Ѐ�?��Q���?��-�7�?O�t�N>�?�����`�?TBP����?J���h�?
ףp=
@|n�b���?B(w}1�?p�j:�?�ⷆX��?�H1�_��?���(\�@��I����?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?<�	��-�?�U'�*6�?4�(�e�?�>���?֣p=
�	@|`�"���?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?�e�:�	�?Dy�5��?��:cc�?�b�X,�?
ףp=
@�j��s��?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?W��#�^�?��I��?      �?	)�L��?ڟ�!T�?��G�z����8I;�?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?����S�?�N�u.�?�&$a��?���7�?      @6�� ��?48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@��j>��?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�����?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?e�Y���?(������?�[����?������?��Q���?{�Z�˹�?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�M���?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?:��]��?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?-����?ӟ���?���;<�?�׷0���?�Q����?���e���?�qV��?�z�G��?�	ϻ���?J��I���?�G�z @��w��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?lt�&��?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?��F�#�?Λ��e.�?�{a���?�D1[�U�?Z��Y���?�z�G�@��V��M�?L�Q���?����S��? 0 ��?4և����?433333�?�a����?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?����g�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�Y��.�?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?���p9�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?�����?IM0��>�?��I��?�h�k��? R���ѿ��B+���?��M1��?�%�8k��?�C���?�������?P���(\�?~Dk���?Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿ���?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?KY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(�w�cK��?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?^e�NF��?�}�K�`�?GT��a�?&Դ���?P���(\�?iS�}s��?����8��?��*H�?>���h�?�؊���?$\���(�?X��WI�?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?gDAl���?<e�U!�?��-��?'u_[�?�Q����?"�R[WD�?�צ����?3�*�" @�#�p�j�?V�;^l	�?(\���(��9���r`�?������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z���c���?y��RE�?n,�Ra�?�$\Z�?��S�p�?�������?��p�4[�?�o��5�?O�o���?�7��ֲ�?J"���?�(\���@������?�d����?���-���?_l�9��?L��N���?P���Q�?�ON���?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�	ږ@��?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�6jDRf7�?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?�'���?�*H^�?�����?Oozӛ��?,\���(�?��x~q��?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?�Gq���?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��?�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?O|-Ϯ��?�SR�&�?}�K`]�?��<d��?w�C�v�?���Q�ο�*UۄP�?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�s����?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�X�!)b�?��h�D��?��P��9�?�1$0��?}��O���?833333�?&~��.w�?T�.�n��?�-�׮�?H{����?������?P���Q�?��/>�?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?���6���?�w���?zkfkl��?�k(���?      @�q�^��?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?��]���?[�[�@�{�q�?.q����?���Q��?�@����? Jx5��?�a�a�?�;x��<�?�������?�Q���@8)���>�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?�S�����?���NV��?��=��?^���?��Q�@�D�y*��?q�l܋��?�������?���k�?t3Q4�*�?�<L�8��?���x�p�?�B-�O��?��Π��?Ȅ�w���?-�؝,��?\\R�M9�?�L8���?=��V���?GҺ���?����t�?�a}w���?H�{�3�?�!>��l�?��m
�?�2�C���?�r����?�M�b�/�?zH��'�? ��(P9�?�&�����?�o$�WW�?��u0(~�?,�x��@�?���\���?񦍺u.�?��?KS��?�Μ�?�� ����?�������?�ۯ<�?
Xl6"��?�Nu~޹�?�
C����?�����Q�?�i2g#��?"���.8�?r��C.�?�*����?< *�"U�?r��E��?��u"��?/���a¿��H��P�?�dRȳ�?�H���?���SU��?�¾���?�Hp:�CĿp�d�y�?���?PÝr���?�֤�Xs�?�;sRA��?Z��TY�?�=[6�?c�w����?`��S�?�п$�?�V|.���?}�����?A��zL��?v �F�-�?�LR�y��?nĞ=:'�?��s��s�?��C+��?9�vș�?`!�F�?�Y��?DX��rA�?6�(���?��|�ѫ�?;�1�x�?Ys�yR-�?��r�1S�?�K�[?��?\�Z���?������?��/��?1%D��?>%����?�/�Bm�?XW�����?<)�Y�?�e��F\�?�<�)>�?���g�?��н<�?�j���?��G��?��-/�{�?�*�x���?/�#�^�?՞���?�����?N.��?��ʓ��?�]��)n�?.�f��~�?�ө�V�?`���[�?2] �?Gz��k�?�RɝV�?ڂ\�3�?�܉���?��s��]�? ���H1�?���٧��?�C�p���?�\dP y�?�H�V���?�~�8r��?ܽ;i 7�?�k�OQ��?T��Ũ �?����7�?��É���?~�Na>v�?(�.c���?���?�;��?"L�� @M�.!��?o���q�?vR�ў�?'&6ꌏ�?�=P�,!�?T�רa�?M�t�d��?{j7��?t
�jR �?l�A����?'�gM�?(�z
�0�?T=���?^2��i�?"�5v\��?B�r}���?Yr�@K�?���w)�?�;Q	��?��z��n�?�g@H ��?��vl���?*�;b�?�� ���?t��>Lg�?=1�Xӊ�?3���?gL�1��?!~��̶�?A���U�?H)�k�]�?l�Y���?��E>�d�?'R��T��? ��A�?����,�?�������?m�g��R�?��@�;��?��봆��?	��2ظ�?EM�BC�?oI��i��?o��	p�?�(6�g��?��g�g/�?(�>���?�Y�-�!�?HMN<c��?E?D[�?%_����?��Y�U�?�A���?�Q�fpO�?���xW��?b׶��?bu�{��?P� &���?Y�b����?�z�#w��?���F�L�?�,'��?�c�]�?�R���?~�|���?t (]�P�?޸N��~�?�vFBc�?��F[��?�B�q	1�?�ُ	k�?/�w*�?`��L�?:�`�"��?��
���?Civ����?S�����?������?�_��k�?��O����?���T�?}�i�T�?F��,�? 2�!��?C������?Z
,�H�?���CT��? ���L�?@t�PH��?_��J��?����U�?�K�=���?�Ĭt~�?w�����?��0ʙ��?�Y@'���?m�3��?�lm���?���{C�?}1A;�?3�zE�?��0t��?��`S� �?y3)g���?K���?��߁f�?1�Rƈ�?�l�us�?�+Et�?����J�?�d�D��?��F(+�?�����?W����?1�ȏ"��?F�hG}'�?��U��.�?�2���!�?�{\���?��s ���?��M�?�	3���?��r�
�?�ۃ*��?�c_ђ�?�GI�[	�?Lnuj�?���d�?�+R��N�?s�,^�?<.Gi���?��h��?�!=!��?x� W�k�?���%�%�?�*�_r�?�R�T���?�͂!j�?��@���?+/���?$���2�?"}{�|�?k�$Ѧ��?��Ű�7�?x~�r��?R��fn�?K7���?�b1o�?�?Tzv/u��?�2�0/O�?��v���?=�U�~|�?��,�Y{�?�XU����?Y�UC�?����{�?Y�[��4�?��yʢ6�?�@�(�?i2}��?�Ceq�?ү4")��?r���ra�?m��i��?�p�He?�v}�5��?��k$�?�_��ؐ�?O�ߔ��?��)��?wAm�ɿY���?½j�r'�?�RU4��?*b(R�[�?nt���l�?Jd�g��?`-��w�?�?�ޞu�?��)Ɋ��?�P� *�?��?Or
�?���q�?]:�b��?�?��HP�?�<qL�J�?8��bO�?���c�Y�?H���ϝ�?��ɶ,�?Q0�][�?�V�e�3�?<� �ID�?y���B�?: ��^��?�)�����?�}����?,�!̶[�? �h3��?��.�b��?
��e�?,�7Ŕ5�?���~2�?G�\"}?�?
u��k�?8�E\W��?�Vk(��?$�Aì��?y�5�(�?��#�4��?�$T�[�?Mw~��l�?
R�$B��?X���v�?3�@o���?��y��f�?�[I�Q�?Z�|���?�G�z�?8��Y]^�?�<�["��?��r�}R�?Oڇ)U�?@0��u��?�G�z�?���;�?�n�3 �?�N�����?�#R��?�� nh��?��69�8�?��(���?	F�r�N�?�Q�C�?��`����?Z>ܭ�p�?��7�r��?p��vp�?��n_�[�?�ylt��?C�ǣ�\�?�|����?0���[��?��<�s+�?ԤH �=�?�Tެ���?�O����?�]��i�?����$@�E�L ��?E�P5G�?~u���E�?�9�xR�?���6��?j�Y2Y�@�p����?�s<�=�?������? .5T���?�X9��?�,;��@X���3��?��ZJ�@�?BtL�O6�?��gh���?Vi'���?r�!|��@�"%��?(�BO��?�ӻ�Fa�?�dĿ���?�����k�?N��@�*�o��?�x���b�?R�GW��?/�VnX��?\^ VaG�?�%>?/N@�UW��S�?��R�H�?n'Z~���?�[w�س�?ZǨ��`�?A��w�c@𵕔��?�$f��%�?�* e�d�?���ꟲ�?E�H��?5�yQ@���2�?�V}��I�?���9��?R���%��?�[�n<�?��}�;@�z��?И�u�?"��+��?�9|(_��?�\N�7�?4�N���?�$2�^��?�:�� �?-�@҉��?�G��6��?vx�.��?���i'�?� IG|�?�Sg}j��?-n��R��?����?�I��+�?P���Q�?d#�u��?&G>7l�?7�2	w�?2��K2��?76���?߬�'��?� �x��?��ݵ��?�������?���jMy�?�l	�0{�?������?����N;�?#d��$�? �&��-�?�8̠��?)�޲�?�j��O�?�����?冞��?�n��i��?Y��/�?Y��X�?�wPNR��?�%���?�s����?�����?s�и���?f�L@���?uh&�W1�?���'��?�?S��?q�eI5�?��4�d{�?,~�Ṭ�?��8)�_����L�Y�?g^+	�?"H>�
�?�_R̆�?��$Y���?�Y�>�?ND��p�?�"�Jի�?p���[��?����?��?%��U3�?�#랅qο�yu���?���
i�?%���-v�?HVk�>�?�T��n$�?F�s7��?�D�!�
�?�ti�s
�?&F(.�?��17S�?��u"�?�Cž�S�?������?C
�ՠn�?��%To6�?þ�]u)�?����E��?i�Q��B�?Ȉ�v���?��K�f[�?r�~,�?Z�9���?����{��?#@�%{��?��O�`�?8��#�? ৣkl�?��ʼkz�?WiE���?)0	X��?rd��n��?< u��O�?b�{[Aa�?P"�J�?��q��?�/E\��?�&�`���?���g��?�*�o"��?d���*��?4��Ie�?�K�^�?�����?/�仮��?'�QE��?����%��?��o��?�WIA3��?�O� ��?b(�ɴ��?���r��?��o[���?r��L4?�?<R/��?hQf[N�?_7dN���?�$V���?ld�3Z��?ad`�q�?��L�D��?�l(_��?6�$
t��?�s���?8N���? �R���?���3�?��� ׬�?^Z���J�?F�d8Z�?�'پ�i�?�w��r�?����@��6�?x�)�W�?���s���?J�u���?�x<�?�o�X.@��ث�F�?#�9Ѕ��?tT>���?�/�	k"�?�|҇/��?$ky�@��.���?IŅ��?1(�;�?���|҄�?=��1^��?�Yĵ�?AFdi��?16����?�ӹ(I�?��괚��?)�lR �?�g����?/[*��_�?�(�"��? �8��x�?���O�w�?I:6h��?i���3�?ʪ���?�,�+ش�?dL�$��?ṋ��w�?E��#��?R��(��?�7���?s�����?3�o�p�?m�t�F��?.�]w�\�?�C��ob�?H�����?b���?��1�S&�??d�$e��?��U
U
�?��Z��?�#�i�?��6���?aL��a�?�����;�?�BP�?p3��=#�?��B��?�'����?�3tfʦ�?X�x���?�����?���Į�?jb����?)�8�Y��?�+=ݗ�?~�菞r�?���'�?�@>c��?���ڳ/�?�#�9���?^�O1P�?�2%�f�?r��g� �?�� 0�^�?�����(�?	ɴ����?Ay����?x�y��?[U�3��?����!�?��"�?��?<P���?�܋=,X�?:{}�]]�?L,qL��?��_�(d�?5��kK�?�_���?�������?�59��M�?�*����?m�r��'�?@>0<#�?�y
���?�06�f�?�Dl�}n�?Cl��K�?�������?_�� �?���K޿�?�����u�?�}Ӈ`�?{�.����?P06Jdp�?s-���S�?u�����?� ��}��?'zk ��?�\o����?	,i`��?��2�S��?<�(��?����r�?Ӡ*��z�?�~�au��?b��b	�?��7����?��Y��?��d����?h�[���?hvZ�8�??F�S.��?�f��_�?������?�=}A�?�duT���?2fs���?�!։�t�?rp�e�?\��I�?�poj<�?�4;.Ϧ�?&��;�?�4�2�n@�E�G]��?]M��o�?;���?%�6I���?�<�64�?���^2�@���\���?���9H��?4-���?�
��Z�?�M�nW�?zo+G�?��]��?����;��?�~�5:��?�T�7^�?�eӢf�?p�i�nJ�?��Җʟ�?�=*����?�|���9�?,��A�@�?�%-�!�?�]�v�?j-�H�?�z�<:
�?�d,�!Z�?�>@��]�?M��jh�??R�+-��?W}�����?BѦ E�??$G��b�?�g�`Z�?/)���p�?@w+���?/�5Ղ[�?�����?�^���T�?fh7�}�?�"���4�?��
A�!�?"���|�?fKŕ���?�Je�H�?_�j��?�I�m���?1]{]�ʿ��߳���?���ݞ�?��m���?|��y]?�?�H#��)�?=�I��̿ï�x�?ʙ8��#�?��S����?�CL=��?�lk��?y�G�ȿ�f���?x�����?�������?>�J�qO�?���%�7�?�D�+T칿6��+eL�?��d���?��Ш~��?�S6�*\�?�����?;��Rӿ{CX�?�ۏ	��?�@jI�?�T!�[��?���V4E�?����#V@4���~
�?қ�qƍ�?���%�?��ޟ~�??MDsH~�?rq#a��@p��@��?5��=lx�?�����?�F�5o�?`<1*��?A�6+�R@�����?m{���O�?��hv6��?����s�?�77ۨ�?��:A@������?JC�_$2�?�������?��t���?�BU���?f�Ѵ��@+|E%*�?�6o�m�?h��P��?\��r��?��n��D�?��3�q@�Zrų�?��#UK�?*�a��L�?b�j���?Y0;P��?�ޮ���@$����?}�u�?t'��G�?�����?�י���?1�Yd�@B$$1��?|� ,=�?cWu���?�l����?
�	*��?�e"�@q|�����?���@�?z%��[}�?7\RYZ��?Z	4��?���E��@^'yUr��?o��oR�?�C��&�?W8��H�?�3����?>�2�-@ο<h��?�쮞�B�?K� 8�&�?(*q���?ъU%���?���P}@P��,7��?�(=z3�?n���?��NS��?�-�ǘ��?����֏@��F%�?����&��?Qrs���?��qzK2�?������?�[N���@!��'p�?Gx��W�?-ծ<H�?��45��?�-��*��?���#s�@8d����?�����?\>�F.��?hUiQ��?���?q�?j�%ŝ@J1e�=��?(%�Orf�?�.%<�
�?���Xt�?��׌�}�?l�X;@(2�p�?�����;�?��!J^�?��܍���?@'[DZ��?��!d�@�ڌ;��?��0��9�?D�Da�z�?�ͨe,�?'�6^bd�?+Nh���@X{��9�?pX�7S�?M��-
��?h����?�/�6�?UQ�Wy"�?];��|;�?<!@���?6���[�?��ټ��?-t��9�?)��%Ff�?b�=H�R�?�8N0E��?�˖���?vy����?���[{�?]�b1Z��?\��o���?��A���?(���,4�?�I�����?­c.���?2O;��H�?$�a��y�?�eu�e��?���I���?��-;��?wWQ6�?+���Ft�?�wG�\��?��6� ��?��p��?�Cى��?ک�{���?�/�K�?�|�@ǲ�?T(�5��?X�{J��?�v�D���?^m����?�����?@���?�u�����? �B����?� 8���?	�ʽy��?�Q��`�?�U��Q��?EL���?F@=����?��ƺU��?+���
�?�^F)��?�w����?Qꍲa��?��t�M��?�{����?�j���G�?P���Q�?i��Xѱ�?�88�0�?P�U�%��?���松�?^݉�L�?}l�U�?�n�ꊍ�?�
�L�v�?=2��2�?�]��.�?d�!++q�?΄|%�?�Hy�x�?�O�O��?Ͽ1�Y��?}�����?aծh9��?�l�v�l�?T��8��?Y�bI�y�?�X�=F�?{	Pc�%�?ov�K�8�?����P��?����N�?+P�DM��?���g��?�#���?�>��e��?`z�B%�?{�=ԓ�?��͙K�?�������?��־[6�?Q�Jj.��?!�>j���?3xT���?��覇z�?a����W�?A���5�?��S���?-��y=��?`A�x&�?��&F"��?>kN']�?�d���'�?�)u�g��?��?�@9��̳��?�-<b��?���r#�?�1���?શwg.�?����6�@��,@e�?�A M9��?�E9x_��?�9�S:��?n7"+��?�Wa�N@�Xx� �?�&�@���?dnV�C��?UG�C��?�����?ڎ�h�@Jæ����?h&w��?/��̈��?�k΂�?��OX6}�?�\l	��@F9���?g��N���?��4:��?$*2���?-��ɣ�?'
��@�� ����?�OP����?Df�n��?X�4l�?��;患�?.�Η�g�?h|�,�?����v��?N��Q�?�`�(��?������?%O��m�?��m�>�?�Q�s��?�&F����?h�R��?�]gs�?��~j��?V{���?l��.���?ƭ�OV�?�H}{>x�?P��/f��?*\���(�?��%���?��4���?��| X!�?���J|;�?k��"uq�?M.�+q�?��ec��?XʾG�?�%쪡1@�ho�?���1�?�<���?������?g�7�?�5����?͖9F�d�?f��@N�?+Bv��?�P�����?������?�Κ�x5�?��B�g�?A� HR@�?�����?��7" ��?�Ny�|��?���Y"s @�@tx���?�������?�OOU���?���5��?�%g�?>%*L���?adW �I�?��-f��?��)y'�?���=��?v&@Ǯ�?0ڧ�Oa�?kvR��e�?����[I�?���D�?�RU�=��?�c_����?�@jw�@4�e$�y�?���(�?�ɤ>��?���l���?ԯ;��?f�K_`H�?^QHn;�?2��K���?1�ȧ]��? (	��?
�Zb&��?B�@0��??�����?!�>E�?K�J�(�@�0�oA6�?�l}����?�岳��?��8�-�?�Zs�R��?x�
'�@4h�6�x�?�m��q�?A���e�?�	��X2�?�%Н"�?~[�֓�@4�K�4��?��*�	��?1l�2N�?�S�E/��? �в�?���G��@��.�9��?J6;��w�? ,B�=|�?�Ng�j'�?��R�:��?�(�>�@1ƙ�7��?9�.�	_�?�9����?#���"�?�����3�?�/�H�?��$�B��?��~�a��?��;|�?2Y���?��J�?�jJ3?��?Ѝ"�qJ�?i4�ۚ�?�S����?%��"��?.o�3��?%š��{�?ν�A��?�	��Q�?"%+��?�o�ϧh�?`�y�R�? ^כ(��?x���?C��3�?a�h#��?!�`�~M�?�z��i`�?��4��?���I��?�͔�[�?��(r�.�?G<�
4��?��S��)�?�\����?�����?A�BQ�?�a����?c<h���?UQ���? Ns����?���,��?�u�M�?��: #��?�?V���?� '[���?�h��r�?��T9�?��0���?"�YZmB�?�Q�����?�>hѐ3�?���w��?Cw�u�h�?��75���?��f�<��?�*,[���?7��N�?��FE+�?�ݭ�k��? 9���?&[L1��?P�����?|�?����?'i�!��?ؘ;��w�?Ѫ�w��?��9t8�?Hq�L���?ٸ-0H��?���5�)�?3 ��{�?��Uq���?"�8(�?ҲN]��?����{D�?M:�#��?#����?�lXg��?+Y���?�Q�1ٶ�?V s7���?lz儁�?"�@q��?���X��?��^+��?W�/��?�jl\�?�$:^@>�?.c�m�o�?YR�1��?`�7��e�?�I�����?(�}����?=�[!�?��eY��?Y�8eY��?̾�\h�?{�vҎ�?��w���?ܻ4ȯ��?J�Ϥ�?�fqU$�?NU����?w+�f��?Eu�w�}�?H�N�@L�D��?��|���?@��-���?��L��?�1O��?w4�-��@�G���?��K`ٛ�?��)�3��?����ۈ�?���:�'�?$@^�i.@/'���?*ӕт��?���M�D�?L�^��?~�b����?�;�US#@�䙗���?:���?b��_�T�?`����?d��\s�?����@i���?- P�	�?��9�D+�?�NH�=��?�W����?Ӣ���z@����k��?�{�WB�?�
ݬ�z�?� �V��?^�����?$g.���?��k-G�?�hj�6�?g����?E:�c}�?�m��.�?�"�Hg�?���t;��?|����3�?rƨ"���?]������?�}ٱ)!�?.(`���?3ӵ�%��?��KcR��?�%hI	 @k���mi�?��Q�
�?R �����n��g�?qEtqFbX
   _n_supportqGhhK �qHh�qIRqJ(KK�qKh<�C�   �   qLtqMbX
   dual_coef_qNhhK �qOh�qPRqQ(KKM��qRh$�B�  !� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _�� d�%���!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��ܶ�pS#��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��Yf�cn��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��b���[���!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _��!� � _����!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@�Ze+�o@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@��!�@qStqTbX
   intercept_qUhhK �qVh�qWRqX(KK�qYh$�C�|�Q��2�qZtq[bX   _probAq\hhK �q]h�q^Rq_(KK�q`h$�CYӃ!Q��qatqbbX   _probBqchhK �qdh�qeRqf(KK�qgh$�C�]�'�ӿqhtqibX   fit_status_qjK X
   shape_fit_qkMK�qlX   _intercept_qmhhK �qnh�qoRqp(KK�qqh$�C�|�Q��2@qrtqsbX   _dual_coef_qthhK �quh�qvRqw(KKM��qxh$�B�  !� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@ d�%��@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@ܶ�pS#�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@Yf�cn�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@b���[��@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@!� � _�@��!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!���Ze+�o���!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!����!��qytqzbX   _sklearn_versionq{X   0.23.1q|ub.