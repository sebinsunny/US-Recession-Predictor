�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?6��C-X   coef0q	G        X   tolq
G?PbM���X   CqK
X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�C!O	� �?qG�w@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?6��C-X   support_q3hhK �q4h�q5Rq6(KM��q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B�                           
                                                         "   $   '   (   *   ,   -   .   /   0   1   3   4   5   6   7   8   9   :   ;   <   =   >   @   B   C   D   E   F   G   I   J   K   L   M   N   O   P   Q   R   T   V   W   X   Y   Z   [   \   ^   _   `   b   c   d   e   f   h   i   j   k   l   m   o   p   q   s   t   u   v   w   x   y   z   {   |   }   ~   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                    
                                       !  "  #  $  %  &  (  )  *  ,  0  1  2  3  5  6  8  9  ;  <  =  >  ?  @  A  B  D  G  H  K  L  M  N  O  P  R  S  T  V  W  X  Y  Z  [  \  ]  ^  _  `  a  b  c  d  f  h  i  j  k  l  m  n  o  p  q  r  s  u  v  w  x  y  z  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                     	  
        	         !   %   +   A   S   U   a   g   n   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �     	      '  +  .  /  4  7  :  F  I  U  g  t  {  }    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KM�K�qBh"�B�K  ���ʦ�?�6f�@��?�~�ϓ�?FM0��>�?�G�z�@F_L�D��?:��8���?�\�]�G�?l�����?������ @�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?s����`�?�0�0�?��e�s��?���]�(�?�������?Eb���?��Y@�H�?�|��X.�?�������?��Q��	@��=�9�?�[��"e�?�+U��R�?�Gq�>�?��Q���?0.Ba��?.�袋.@�
�l�?haz�g�?      �?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?�jǊ��?������?<�7b��?"�r����?أp=
�	@^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?F}�p �?������?N6����?\����?ffffff�?��ԩ/��?AR˔���?JL �F�?�>,��?�������?E��.��?5�\�`��?���nD�?P��n��?�(\���@�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?W����?��8��8�?      �?Au���?�������?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?������?�{�D!�?�l.�VP�?�2��h.�?)\���(@���*�_�?۶m۶m�?E������?�n���?�p=
ף@0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?"K�_y�?���,d�?���<�?jhɬ�?�Q���?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?9�KO���? ���?R-ŭX�?X�,)D�?\���(\@�!K���?)^ ���?u�`6�?���j��?q=
ףp�?^���*�?Z5�Uc[�?���l��?Ҏ#��?�Q���?R�p,C.�?������?��U�	��?n��x�>�?��Q��@lv��?*.�u��?m�����?O�<�"�?!��Q��?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?���#�?})�Z�?d#D:��?��;�?��(\��	@�Fm�}�?�/Rm���?q�Q>	�?ݫ`���?=
ףp=@-����?ӟ���?���;<�?�׷0���?�Q����?Qn�p&�?�؉�؉�?�*����?��M�`�?�p=
ף@��i�,�?ףp=
��?���b��?,Fڱ�?��Q�@�y]>d�?g;>)7�?�Ǭ�NR�?&H-/|�?=
ףp=
@�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?i�+s�?333333�?`�>��R�?��.���?q=
ףp@L�|9��?m���X��?�B�q��?����:.�?833333�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@e�F-��?�������?���:%�?V���g�?ףp=
�?EÓ���?�����?�&z��V�?WUUUU��?���(\�@@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?�t&����?��(��(�?�^mSz��?g�Bg�B�?������@�c��)�?c��4�?�.fxx�?�Ŗ����?������@�Dz�:�?�=��!�?���f�?�%��}'�?�p=
ף@�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?x����v�?4H�4H��?�)~�r��?���Kh�?�p=
ףпm�<�?     �?�������?A�zy3A�?{�G�z
@"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿ���,��?ى�؉��?��� W��?{�G�z�?*\���(@,"�j�%�?,-----�?'狗�8�?�`�����?133333�?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?����-�?��L��L@;K�*�O�?��
��?�������?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?�����?IM0��>�?��I��?�h�k��? R���ѿ/9(��?.�袋.
@�*����?�������?�������?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?Se�;f�?h����@A�j�}��?�WJ�B��?S���Q @��Zb��?��+x���?� �Y]��?����?hfffff@��;�l�?��{����?��`|��?���!�?@\���(̿濸����?r���0�?,�C ^��?5���4�?���(\��?톘��=�?+P�W
��?���gk�?�������?Z���(\�?��y����?I`�:�?�5G��`�?4h��J�?      п�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�ۇA�?��*�3��?���R�]�?AA�?��(\���?Um�����?�t��N��?�;1��?_�1yo|�?r=
ףp@�@��+W�?��)o���?�߾���?      �?������@��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�?�wF�?��D'�?6������?�_�_�?�������?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?���Y�?�	g�	g�?ya��w�?!s��2�?�p=
ף@r6]����?�������?�	��6f�?���3$��?H�z�G@S\�C{��?5�rO#,�?64�����?�|�G�j�?ףp=
�@<�	��-�?�U'�*6�?4�(�e�?�>���?֣p=
�	@��2���?���?��</�b�?�ռY͛�?H�z�G�?48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?��sr��?��3���?�V��?��~5&�? ףp=
׿���?�m۶m�@��X)�O�?�\.�?)\���(�?dwl���?d�fI�m�?��W�6\�?=]�:��?)\���(
@���e��?I��/�?i�(�U�?�VC��?T���Q�?�4��
:�?(6$�)G�?(��J+z�?v��4��?���(\�@�������?�m����?G��|���?E4Z����?�z�G��?W['s�,�?E�JԮD�?��K�y�?��J�[��?r=
ףp@�N"H��?����?Hx`2��?��r:���?������@�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?����?1bĈ�?��6-f�?�Ab�k�?�������?�>����?      �?0`z��Q�?'u_�?�p=
ף�?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?C�Z����?�Nu�w��?��سX��?�R:CW��?H�z�G@�u����?�wK�?��?�ef���?tT����?�z�G��?
��\���?��\AL��?)us�?      �?433333�?���g
�?&���^B@���X^�?��FS���?G�z�G�?��S��?I�$I�$�?�����?���w��?�������?�h�{���?-��K���?滵P�K�?��)W]��?q=
ףp�?
�&af-�??�?��?�q-���?��	�{�?أp=
��?�4~���?h}�}-�?	+��]��?�ܽ*���?�Q���	@�$�vQ�?����?dȇ���?�?2�խ�?*\���(@���� �?�$I�$I@W�G#��?"1ogH��?ffffff�?O@���?ffffff�??w��a�?�A���?��Q���?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?r�2�F�?�zۜ��?z!I�,�?c[:��c�?�p=
ף@
��@��?���Қ�?'::V�e�?��JR�?������	@�Ĭ~��?��Q���?>s=��^�?�����?�(\����?:�X{��?���.{�?P�l�V��?'��,�?      @s��&�?(W�7�?���xW�?B�HV��?��(\���?}��Yc��?���_��?+��6rl�?W�m���?�G�z�	@�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�2�j���?     �?u�;�F�?�$I�$I�?�z�G��?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?b�+d�&�?�L�w�?U�&xl�?=��k�?�(\���
@z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�
>U�?
ŭP�
�?Pf�i���? i]���?�G�z��?:+��?NB�3�?Ci!��?r�q��?Y���(\�?C�oB��?      �??��(b-�?b�1`�?433333@R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿW#Q�.�?贁N�?��W9��?�$A��?!��Q��?��p����?      �?��e�N�?�������?R���Q@K�^�/�?(✭��?.�, �y�?!z|��?R���Q@�4����?�%����?�J:��?v{�e��?���(\��?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?�\7z�?���"��?����}�?7�j�?H�z�G@��9���?�e���?��G��\�?�����\�?���(\��?8����?�gS��=�?�~��H�?�Vi�_�?�������?Z�yv�<�?��a�
��?��ࣹO�?:&߭��?��Q��@��(��?7�Y�"�?ޤ�=%�?{�!���?���Q� @@i���?P��O���?�k�9���?��U�^�?(\���(�?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?aC�����?     �?J�.����?"1ogH��?��(\���?�מ���?�i�i�?Q�XW��?�R�~���?      �?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?(1B���?b'vb'v�?s�ӭ��? �R{���?H�z�G@��_O�?��G��=�?�!|����?L��7���?033333@)��h��?UUUUUU�?�����g�?�X>b��?���Q��?� �9�$�?h���Q��?�3�s�?�B#�E�?��Q�@�}��?       @j��_�?��¯�D�?�(\����?�$�l���?d!Y�B�?k���?"�?d�*|��? ףp=
׿ 3`���?���P��?�D�e'~�?�]���?{�G�z@9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?�p^��m�?tT����? ����?����x�?���(\�
@����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��;4��?WUUUUU�?��J�l�?W�m���?H�z�G@��Ʀz��?��*�{7�?�
���?�o��o��?733333�?'�CU$
�?      �?�t�U�%�?.�#EC�?��Q�@Un����?�������?#�R���?]�����?�Q�����%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�C����?�������?A�ra���?�@۽U��?���Q��?�y�]��?]�)~I��?��@��[�?�{����?���(\�@���~�?9"�P9�?<O�����?!������?���(\��?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?��,���?�z�G��?����U��?a���{�?      �?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@�x�\�?��2����?ؔ�
&w�?      �?أp=
�@�D̥�
�?�Zk����?��iz�?���\��?��Q���?-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?��L��?�q�q�?G`3�!�?O���t:�?R���Q@szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?��X���?l۶m۶�?�r/js�?]t�E]�?���Q� @=��a��?}T$;f)�?�|��O�?�UO���?��(\��@EtA%�?/���}�?�f�M��?��¯�D�?���Q�@%�����?*��RJ)@f|��O�?D0��fa�?�G�z�?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?�m�=���?WUUUU��?���a�?v{�e��?���Q��?��A!K��?r�q��?�=�� �?�١�?�G�z
@����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?��״��?Ѻ���@��O��?����T�?���(\��?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?_^MiK��?�q�q�?P����?@�wܛ+�?\���(\�?)�x�?UUUUUU�?JB��EX�?�-�t�b�?q=
ףp@����?CBq�n�?�M���?ABЋf��?hfffff@=B�k��?g�K1_h�?;9�=-�?$�D"��?q=
ףp�?���|�?      �?��`��?iiiiii�?{�G�z@����Z�?+�O��d�?���s�?���rD��?������@�|��	�?b�־a�?pA�D�?���rȔ�?H�z�G@a�B��?�������?' Z�u�?�����?���Q�@P�����?UUUUUU�?�k�1���?O�n�	�?��Q�@��j�G�?u�5�o��?���d��?�~��?�G�z��?Za�T�
�?�1���N�?D��car�?�MҷV��?H�z�G@:N�1��?G�:y�?Y<�&!�?F����?��(\���?�o�����?��%�̀�?�\"�0�?P[AG:��?�(\����?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@����?      �?ŵ�a��? )O��?      @2�7���?���A�?���i���?_7��T�?R���Q@c&i�?�ÔP��?P>�z��?�uI�ø�?      �?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?\��Z�?�$I�$I�?��ԉ#\�?����>4�?]���(\@\�f��p�?� ���?�Z���?�Ytl�?�G�z��?������?������?�X^o�?��<t/�?H�z�G�?4s���?�����?/z�V�4�?~"����?H�z�G�?���[�?����NB�?b%c�r�?����]�?hfffff@�܎h�?��/�$�?�p\��?���6�?���(\��?�J�LT)�?�������?5�Z(��?XV��?��Q�@�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?ϙΔ�?a#@i��?M��d�?��,��?      �?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?evoƃ��?�q�u�?�)���R�?t������?0\���(�?L�Q���?����S��? 0 ��?4և����?433333�?�l���!�?�9�s��?�1�[x}�?�[��"e�?*\���(
@_i�"�?VUUUU��?��i��?)\���(�?�������?t��!���?,�X��?^*��U��?�:�>c�?��Q��@W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?���S��?��c�0��?k��{<j�?9
�
0�?<
ףp=�?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?����q��?      �?M��7���?      �?�G�z @X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?�
⛏A�?��P���?4 ��<�?(
P�;�?������@��t�j�?��qg	��?d���1�?(�)��;�?�������?�T����?Z7�"�u@m�����?����T�?�������?���1�?��fy��?���N�R�?Wŵ.���?���(\�@���n��?�n0E>�?T3	Z�e�?xH����?R���Q
@�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�W���?{�n��?	sG�h��?в�9��?��(\���?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?[��`��?ك2�*j�?� �;��?�������?�(\����?P,��v�?�������?4:�$�x�?�%����?�G�z�?��*�?9�&oe�?ߘ�[]�?��Я[[�?��(\��@y�-[Y�?�8�?'�8����?%���E�?�G�z�@����?�N̓���?�[����?*) �'�?\���(\	@��I��?      �?	)�L��?ڟ�!T�?��G�z���0k��(�?�Iݗ�V�?���Y&�?���?�?      �?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?T,���?T:�g *�?"�[��t�?7.Hj��?�������??d~-��?�u�����?����2�?� ?7��?      �?E�X9�x�?-��,�?)=��'�?��0���?�Q����?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?{��*W��?     @�E!��p�?�$I�$��?�G�z��?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?�r�>J�?�|���?n1DE-[�?|�,����?�z�G�@@>`]p�?;�;��?�����?���O��?������
@�O�<�?������@uq_�E�?��$2��?H�z�G�?����em�?׊��+��?Y�����?"$�A���?�(\���@�83���?�{Nm{�?�F�� �?�������?P���Q�?��0��?R�}�=�?ӗYl�n�?.�袋.�?�Q���@}v�Ʉ[�?y�5�װ?X/�$R<�?8��Moz�?)\���(@*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?3�J���?�F�tj�?^���i��?�
� ��?�Q����?��=O�?M4�DM�?���2��?�ܛ���?
ףp=
@{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�������?�$I�$I@��;���?R���Q�?�z�G��?N"����?FFFFFF�?�-5��?����o�?��(\��@뀂���?��Bt�?�(�=l�?��ұ�?أp=
�	@Po�S3�?!1ogH��?�8Sn�Z�?8Q�H��?�Q���@!��m#�?r�q��?�_پ%T�?"Y�B�?{�G�z@T-����?UUUUUU�?L�5���?�������?ffffff @@�X兞�?f���?����15�?�>��?��Q���?փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?����0��?�x��ܷ�?Y1"�	l�?l#֥���?��Q��	@�n���?H���x�?6?�x�o�?�#�	<�?R���Q@erV�lw�?�6S���?�q9˲��?%�e�@�?�p=
ף�?�'=��?��fě�?��Xf[�?���¯��?�G�z @6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?Q�����?I�$I�$�?���Y�?z��!y�?333333�?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?�@����?�����?���Q{�?(������?�p=
ף@5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?��� ��?:��8���?��'c��?�-Wr�?333333@�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?��S3;��?ĸ_�T>�?��a8%��?�,�י��?q=
ףp@O�TE���?�(፦@��x�b�?��RJ)��?�������?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?�_����?      @����,��?[�o�W��?���Q��?8P��A��?�\;0��?<b���e�?y{�X�?      �?~�W�f��?y@�z��?�{b�?�W�^�z�?�z�G�@I��q��?�'iq��?�&��?#�����?�Q����?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?0	�`���?o�vu�?N�� V�?��X���?��Q���?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?mӞ��?#��~j��?�1?��l�?��i���?�Q����?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?���RG��?"�u�)��?��s��?��o����?�z�G��?�h�(���?����?�3��=�?g�=���?�������?��zZ �?&jW�v%�?t���?X`��?!��Q��?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?��n9�
�?�Zg_D��?_j�P�?r1Bm��?H�z�G@_�;I*��?k��FX�?e�5���?J����?R���Q@�{����?�Pd����?�{c����?�������?���(\��?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�?;�H�r��?W�rCH�?��A�^�?�����?(\���(�?�]�L�b�?2&�l�?      �?]|�c���?�z�G�@�va�q�?iiiiii@�;��`�?      �?433333�?�G,���?�	����?���R{�?��?�c��?���Q��?G�u���?�t��6�?ZM��W�?�ɵ��?gfffff@{^Q�h�?       @��Tf,�?�7�7�?�G�z @�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?Sª����?      �?�	*�/�?W�<�?R���Q@5~�lk��?u32"��?8����j�?�����?�z�G��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��Sr��?U����?<����?w�{��?<
ףp=�?��aJ��?��˝��?�D�y�?�$���?���(\� @u�-BK�?��T��K�?��x���?>���~��?���Q��?e�Y���?(������?�[����?������?��Q���?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?}9�ot��?d����.�?֐��<�?OP�?�z�G��?%���y��?a8B��?�!!?�Z�?���q6�?<
ףp=�?����*�?)#�`��?��@�x�?�gL���?أp=
�@:����?�5��P�?v$����?;�;��?أp=
��?��]��S�?�z�����?����?1�0��?(\���(�?6%�M���?���s @N�|ҍV�?e�e��?�������?� �����?{ӛ����?��*��I�?"�nd=6�?������@�jS`��?&o7�-�?󇕔p��?N�K�?�Q����?Ũ���?WUUUUU�?%�[P�~�?�������?�(\���@�m�02��?;r����?���	���?����<�?��(\���?"ۼ7@��?�q�q�?=ȋ��?H�z�G�?{�G�z�?�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?����t�?���j?�?��y��X�?sƎ�e�?������@E� �?      �?��ԉj��?��|�nS�?333333	@��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?|A� *��?�袋.�@��k{�?W�+���?H�z�G�?��r���?\��[���?�4�.��?2}~k���?��Q���?��X��?�Kh/��?�f i5�?*g���?���Q��?��1���?wF]�K��?={��?������?�Q����?���X �?�\�\�?6#�|a�?>6:8���?P���Q�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?��;��?*b�����?�0����?�8+?!��?���Q�
@,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?�j�с�?�dn}�?�xJ�Rn�?��寖�?�z�G�@X���A�?������ @<�z^��?C���,�?�������?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?��{G�?����S�?Y�_��?�����B�?֣p=
��?�!ފ�?c����?��J%%�?��(\���?�G�z�?]��{��?�����?Iy���?E�,V!�?�Q���@h��Ƅ��?UUUUUU�?���t�?     ��?q=
ףp@S;>���?�Y���?�gS���?U�j�o�?أp=
��?�����X�?t�����?�^Y�?��??��5���?ףp=
�?P�H �?:��8���?Ta�z`�?�'�����?�G�z�@�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?əPB�?��.���?gL0�h�?l��(�?ףp=
�?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?V�gb�?��W�l��?U�����?_�HI��?�������?��/����?���T4�?h�v�Q�?�����? ףp=
����B~���?ƶ#e��?-��k4�??&ǒ::�?{�G�z@ '�Q�^�?ᖚ�?C�7�y�?4H�4H��?���(\�@(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��<���?      �?��(�r�?��a	G��?���(\�@��m��?����?&z`�5�?2u�=�S�?      �?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?
��Y0�?�G*;�?      �?������?��Q��?"&�H
�?�?�4��yO�?��)��?
ףp=
�?/������?�k��%�?���g���?8S����?�G�z���0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?~�aE�?"�z\��?�R����?I��/�?.\���(�?ӏK�K�?��{���?���S��?{���g�?P���Q�?wJ��L��?S��?�p���?�������?
ףp=
@�X��S��?      �?Ѹ�U�?1�0��?���Q��������?�Qf�,�?z�<���?�%���x�?Z���(\@r>bܘ�?��MmjS�?e�����?|1����?���(\��?q�ک��?      @���<X�?��=���?333333�?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?�uf�K��?EDDDDD�?ޮ@l�Q�?�������?      @n,���$�?����b)�?A�쎑��?@�1���?
ףp=
@����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?�_�^�/�?      �?K��>�?0�9�a�?������@P@��}�?��k���?      �?�J���?�������?Λ��e.�?�{a���?�D1[�U�?Z��Y���?�z�G�@�miV���?�U�;���?P�l�V��?A�Iݗ�?�z�G�@뚖f�?1ܫ`���?��Z(~�?�;�;�?@\���(̿Y/�7�/�?�>�J�?��	���?t�����?���Q�@���]�?��g����?1sJJ��?��f$/��?���Q�@�]A6�?��0�:�?A�B)���?7��O	�?�G�z@�����?�DxR���?`f�"�?�8yh=�?q=
ףp�?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?*����?{���\�?�N�ҝ�?�����?�Q���	@XD"���?R��+Q�?$ ����?�#F���?P���Q@��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?����g��?�]����?P�øW�?v�=H]��?��Q���?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?auȒ���?�v%jW�@��s5��?`����?�Q����?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?�74J�_�?*6\u��?�$8����?�/t���?      @����?���a���?Û�P�?�`8wC�?P���Q�?�p�|���?���)��?^�3���?h�J� :�?�Q����?l,����?gH���?���2G�?v�A����?�z�G��?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?����?��R�y�?�����?�s@ڦ�?�p=
ף�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?������?�~H���?U��oW�?��S�r
�?
ףp=
�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?������?�5��P^�?lN�b�Y�?���v�?�G�z�@D���Oz�?PuPu�?      �?٫��J�?���Q��?������?�N��N��?��U>R
�?	f���?�G�z@T�.�n��?�-�׮�?H{����?������?P���Q�?�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?*�fV=�?'���?<��v��?ZLg1���?�������?����8��?��*H�?>���h�?�؊���?$\���(�?�����?)�����?�s�H�?�u�y��?�G�z�?�r*��?z�Ha��?��R����?�{mĺ��?���Q��U@�'��?�x+�R�??dM2_�?�(S�\��?�(\�����п�cX�?���؜��?��{�z��?�F��?_fffff�??V�)��?_�_��?      �?��B�
�?�G�z�?¶�F�s�?0w�fs�?)���k�?y�!���?{�G�z@\�����?�3�u�?�d�yv6�?f����?���(\�ҿR8�u�?S{���?��,�1�?:�oO�$�? �G�z���qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?(� .b��?�k�S��?��F����?���w���? �G�z�?fo/���?/����?'N`�4��?��3���?�����������C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?��bK��?�/��/��?T��cP��?.Ԝ��?�Q����?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?Ե7�rL�?�l��l��?���'��?��E���?��G�z��g�\���?�����?��񍔎�?����.��?�G�z�?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?���6���?�w���?zkfkl��?�k(���?      @�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿:M�]��?HA@s}�?g0�d��?��7���?\���(\@�X$����?L�:,��?&����?G�N��?\���(�?I)i���?�{0�I��?KU���?�X�����?@
ףp=��i����?T����|�?�;x�]z�?,d!Y��?P���Q�?��h�D��?��P��9�?�1$0��?}��O���?833333�?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?y��RE�?n,�Ra�?�$\Z�?��S�p�?�������? �	�'��?pN�F��?�^mSz��?�]�P�?�(\����@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?+e��R�?pА����?�_P�
�?���譺�?��(\���h�����?��1����?�IF��?�_{�e��?��G�zĿ�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=�KY,i�a�?�$I�$I@2�ܫ���?OV��ȫ�?(\���(�������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z��G���;�?�x+�R�?gj��?�r4.G��?��Q�@�ao�2 �?�Λ�~b�?����?H݊ÿ�?���(\�ҿ(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?�ݭ����?yþ�\�?�CM`��?�w��K�?�p=
��?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�'���?�*H^�?�����?Oozӛ��?,\���(�?�S�����?���NV��?��=��?^���?��Q�@�o��5�?O�o���?�7��ֲ�?J"���?�(\���@�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?Mt�å�?�k���?#�%%ֆ�?�u�)�Y�?������ɿlq�����?ѭ8��7�?�V8Y+��?��07�Z�?������ܿ��K���?8F�ʹ��?�U�K���?��k���?x�G�z�?�d����?���-���?_l�9��?L��N���?P���Q�?P��-��?�NV�#�?8��m���?�;�#�?333333@�q� .�?��"E��?�V���2�?�^�^�?�G�z�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?��]���?[�[�@�{�q�?.q����?���Q��? ��2�?S�n0�?���&�_�?I%�e��?�������?� �����?r�q��?܌��! �?���[���?��Q��ۿ�깘4��?�7M�?�i�'��?$p�?b�?=
ףp���[�à�?��b����?��y�xi�?�cp>��?�z�G��?�,��o*�?���tT�?Eg���?�@i�
�?���������L���z�?X�O���?��F�{�?!���c��?�(\����?[�_�?r���&T�?Vl;!t��?�O��O��?�Q���?u��=M	�?�ڧΪu�?f>����?: 2ܫ`�?�p=
ף�?v��� �?o}$�o<�?��(ET��?�{i�"8�?���Q�
@����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�`���`��?���-��?����w�?��-�jL�?��(\��ſ��B\&�?�n0E>��?���L�?2 K��?�(\����?[̽e��?�)`>�]�?i���/��?o��[�?������?���fR�?:�:��?�Pk����?ק�����?��Q�	@�+����?�#�;��?��oa��?��8���?�Q���ѿ_������?���h��?�����?\t�E]�?�������?F��W~�?��f=Q��?�����?DDDDDD�?P���Q�?��
�?�"nps�?�`>J�?/������?���(\�ҿqCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�  O   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM��qPh"�B   颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���0�y����颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���颋.���fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@fMYS֔>@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�C@]����y?qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�C�ŭ6�`�q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�Cc��m����qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�C@]����y�qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM��qvh"�B   颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@0�y����?颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@颋.��@fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�fMYS֔>�qwtqxbX   _sklearn_versionqyX   0.21.3qzub.