�csklearn.svm.classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX   kernelqX   rbfqX   degreeqKX   gammaqG?6��C-X   coef0q	G        X   tolq
G?PbM���X   CqKX   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   f8q K K�q!Rq"(KX   <q#NNNJ����J����K tq$b�CX驅���?�S�n@q%tq&bX   classes_q'hhK �q(h�q)Rq*(KK�q+hX   i8q,K K�q-Rq.(Kh#NNNJ����J����K tq/b�C               q0tq1bX   _gammaq2G?6��C-X   support_q3hhK �q4h�q5Rq6(KM�q7hX   i4q8K K�q9Rq:(Kh#NNNJ����J����K tq;b�B8                           	   
                                                   !   #   $   %   &   '   (   )   *   +   ,   -   .   /   0   1   2   4   5   6   7   8   9   :   ;   <   =   >   ?   @   B   C   D   E   F   G   H   K   L   M   N   O   P   Q   R   S   T   U   V   W   X   Y   [   \   ]   ^   _   `   a   b   d   e   f   g   h   j   k   l   m   n   p   q   r   s   t   w   x   y   {   }   ~      �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                 	  
                                   !  "  #  $  %  &  '  (  )  *  +  ,  -  .  /  0  1  3  5  6  8  :  ;  <  >  ?  A  B  C  D  F  G  H  I  K  L  M  N  O  P  Q  S  T  U  V  W  Y  Z  [  \  ]  ^  _  `  a  b  c  d  e  f  g  h  i  j  k  l  m  o  p  q  s  t  u  v  w  x  y  z  {  }    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                   
                              "   3   A   I   J   Z   c   i   o   u   v   z   |   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �                    2  4  7  9  =  @  E  J  R  X  n  r  |  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �    	  q<tq=bX   support_vectors_q>hhK �q?h�q@RqA(KMK�qBh"�B�b  �v���?U�����?����?�M����?�(\����?2�g2��?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?I)i���?�{0�I��?KU���?�X�����?@
ףp=������?����r3�?Q@����?�.���t�?A~�9�J�?�p=
ף
@I��~0�?�r��Φ�?�n�l�N�?0��x��?3m���G�?|�G�z @�du��x�?w���2��?Z7�"�u�?D����?�h�Q�&�?8
ףp=�?8K����?m��C�?      �?2zW�]6�?��L��?���(\�@��y����?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?�i����?T����|�?�;x�]z�?,d!Y��?P���Q�?���}�I�?~�aE�?"�z\��?�R����?I��/�?.\���(�?�&�s�n�?Q�ps[-�?#N�	���?�[�����?��)��
�?������@@� �,�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?�0�P��?c(x'�?�l.��?!YY��?�G�z�@|�0l+u�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�9��-c�?�j���?�B��X��?�����0�?.ܴE�?��Q�@Ec{�'�?�m�=���?WUUUU��?���a�?v{�e��?���Q��?������?-B�h�Z�?�$I�$I�?���_��?��|��?\���(\�?v�����?��mW(��?333333�?"�*|��?���?333333@��K���?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?H��O �?���C��?£^b֑�?���;�L�?�z�G�@6ۮܹ��?J��:���?=
ףp=@��=!E�?���E�?=
ףp=�?O����?��39�??�?��?��¨���?;�/,��?��Q�@�����?_^MiK��?�q�q�?P����?@�wܛ+�?\���(\�?ǘ8�+�?n#�{�?%z�$z��?0�1��k�?��M�<��?      @Zvr7�6�?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?
��\���?��\AL��?)us�?      �?433333�?@�����?\��Rx�?�ۚ��?�<�}C�?����C�?H�z�G@H������?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��? �	�'��?pN�F��?�^mSz��?�]�P�?�(\���近x����?^���O�?o��o��@�H<�'�?�X�%��?�������?�8�T/�?����?���a���?Û�P�?�`8wC�?P���Q�?���Z���?��y����?I`�:�?�5G��`�?4h��J�?      п�P�$��?���*�_�?۶m۶m�?E������?�n���?�p=
ף@�CUK��?փ���?�L�w�?���tA��?��pHJ'�?@
ףp=�?����y�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?t� %��?.�袋.�?����2`�?��H	9�?=
ףp=@�ө}���?S\�C{��?5�rO#,�?64�����?�|�G�j�?ףp=
�@ �K.R�?��n9�
�?�Zg_D��?_j�P�?r1Bm��?H�z�G@,2F:��?Y/�7�/�?�>�J�?��	���?t�����?���Q�@8�ϵ�/�?%�����?*��RJ)@f|��O�?D0��fa�?�G�z�?����խ�?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?y�N�?�'��m�?=J�i�?     8�?      @v�u����?��X���?l۶m۶�?�r/js�?]t�E]�?���Q� @�XJ�N��?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?����g�?����?�N̓���?�[����?*) �'�?\���(\	@]�l����?R8�u�?S{���?��,�1�?:�oO�$�? �G�z��S�hz���?������?�~H���?U��oW�?��S�r
�?
ףp=
�?���y[�?8����?�gS��=�?�~��H�?�Vi�_�?�������?�11�G��?<�	��-�?�U'�*6�?4�(�e�?�>���?֣p=
�	@|`�"���?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�)2��W�?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?:r����?��S��?I�$I�$�?�����?���w��?�������?ݝo��?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?����Z�?r��Z�@� ��r�?g��|�Q�?033333�. }0�b�?O�t�N>�?�����`�?TBP����?J���h�?
ףp=
@|n�b���?���`�?��`Q�(�?w
R�VO�?�>���?)\���(@���я�?�\7z�?���"��?����}�?7�j�?H�z�G@�N���K�?�aݚ
�?(������?� R�M�?��7��M�?       @St��i��?��8�N�?�L�w�?4��z��?i ��[��?�p=
ף
@�M**ˋ�?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?�@�,��?I�$I�$�?x�?q�?u<@�La�?\���(\�?�?i���?����0��?�x��ܷ�?Y1"�	l�?l#֥���?��Q��	@S[~f�?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?���|7�?ۍ}��	�?>}���?��ũq�?��������?:��z�?�p�|���?���)��?^�3���?h�J� :�?�Q����?���ah��?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?��p����?      �?��e�N�?�������?R���Q@>����?������?�ߥ�l��?��7v�?�c+����?q=
ףp�?����o�?֊�q��?��Z��Z@�K��?#e�����?���Q��?
k#w��?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?*��Al��?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�?�p^��m�?tT����? ����?����x�?���(\�
@:�%�?*����?{���\�?�N�ҝ�?�����?�Q���	@WV��u�?J��YL�?VUUUUU�?!��a���?�7�7�7�?      @%CE����?���%�?������??�0Yp�?��ퟡz�?r=
ףp�?Y��γ�?��S3;��?ĸ_�T>�?��a8%��?�,�י��?q=
ףp@p��8�?Ũ���?WUUUUU�?%�[P�~�?�������?�(\���@4���x=�?e�Y���?(������?�[����?������?��Q���?{�Z�˹�?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?Ψճa�?j�^�c�?���2�?cA^	}6�?أp=
�@���ي�?\��Z�?�$I�$I�?��ԉ#\�?����>4�?]���(\@�6L5M�?�ꍑ��?�h�����?Xn�e�w�?��:X���?�G�z�@���{��?����?      �?ŵ�a��? )O��?      @�����?evoƃ��?�q�u�?�)���R�?t������?0\���(�?I��p��?��E4�?Dio����?J_��_�?�����?      @�ۚ%+��?�ӄ���?R���Q@���K���?����*��?�(\����?I^J��?O@���?ffffff�??w��a�?�A���?��Q���?j�úg�?wJ��L��?S��?�p���?�������?
ףp=
@�9e���?"�FU��?�71}�?v��3���?�N�Q�S�?�Q����?�5�,[�?���E�]�?WUUUUU�?��o3��?p-ܴ�?��Q��@h�:� ��?`���`��?���-��?����w�?��-�jL�?��(\��ſ�E]�?�����V�?6����?�xf��??�����?������@C2h�O�?�+����?�#�;��?��oa��?��8���?�Q���ѿH����?��9���?�e���?��G��\�?�����\�?���(\��?:����?�$�vQ�?����?dȇ���?�?2�խ�?*\���(@��W���?��t�j�?��qg	��?d���1�?(�)��;�?�������?�O^J��?P,��v�?�������?4:�$�x�?�%����?�G�z�?Qj����?!��m#�?r�q��?�_پ%T�?"Y�B�?{�G�z@����?���Y�?�	g�	g�?ya��w�?!s��2�?�p=
ף@n�5��?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?�=�,;��?!G%޸��?������?ُ�؏��?�G�z�@������?@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?i�o��?oCӱ�>�?Y�eY�e�?�}{�:��?�p'�p'�?������@�?�����?��=Qr�?7r#7r#�?y�sJiM�? ��c��?433333�?�Qa���?�@����?�����?���Q{�?(������?�p=
ף@4��6I�?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?���A��?m�<�?     �?�������?A�zy3A�?{�G�z
@@s���#�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?�徦�<�?�\AL� �?      �?�������?��Q��?�A���?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?�D�;$�?���&�?�p߃���?��N�M�?�G�z@ԫ�|$�?��aJ��?��˝��?�D�y�?�$���?���(\� @��p��A�?� �����?r�q��?܌��! �?���[���?��Q��ۿ�#Bt�?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�b=��
�?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?���S��?��c�0��?k��{<j�?9
�
0�?<
ףp=�?z��w
�?�uf�K��?EDDDDD�?ޮ@l�Q�?�������?      @��E�E�?2E�Ĵ�?	��-��?'m�`�?:o1���?hfffff�?��E T�?����?��Pp%��?kub�Q�?̟�Ѐ%�?���������X5�Q�?&�-ʰ�?�.]�6�?���}���?K��0a]�?������@�MU�Ǖ�?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?��L�F��?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���?g�\���?�����?��񍔎�?����.��?�G�z�?'�����?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�`1+�H�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?�9ɻ�	�?     �?vc���?�;�Y�?q=
ףp�?�e���C�?F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿr���;�?����t�?���j?�?��y��X�?sƎ�e�?������@~��CР�?�����?�Qf�,�?z�<���?�%���x�?Z���(\@��w]�f�?P5��3*�?Y�eY�e�?/�G�a�?�M6�d��?H�z�G@I��sR�?��{�A�?,˲,˲@�Z�rf�?c��0u��?���Q��?��v��?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?Za�T�
�?�1���N�?D��car�?�MҷV��?H�z�G@Ƨ�/5��?�*�N��?
ףp=
�?_�6�?:����R�?�p=
ף@}�"�>�?���X �?�\�\�?6#�|a�?>6:8���?P���Q�?��f���?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?|? ��@�?¶�F�s�?0w�fs�?)���k�?y�!���?{�G�z@��VFr�?��[y��?�Ў�e��?��^*)�?z^{�?�(\����?�9)�?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?�H�9���?�oX����?�%oV���?�Fn�Fn�?��Q��@�m�J�%�?�Ĭ~��?��Q���?>s=��^�?�����?�(\����?�a��~�?C�oB��?      �??��(b-�?b�1`�?433333@��
�f�?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?u��׿�?U[G[��?;�;��?�	v�o�?�a�a�?������@U��A��?�S�����?8�P\�?��;^�?M�*g��?\���(\�?�	�;D�?����-�?��L��L@;K�*�O�?��
��?�������?��R{~��?����em�?׊��+��?Y�����?"$�A���?�(\���@K������?Λ��e.�?�{a���?�D1[�U�?Z��Y���?�z�G�@��V��M�?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?�miV���?�U�;���?P�l�V��?A�Iݗ�?�z�G�@خ�V��?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?g?�V.�?z&�����?�H(m���?��K�y�?���cY��?��Q���?��ʦ���?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?{��*W��?     @�E!��p�?�$I�$��?�G�z��?�_�����?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿|�TT�+�?ӏK�K�?��{���?���S��?{���g�?P���Q�?�Z(O,k�?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�??[�w(�?� �����?{ӛ����?��*��I�?"�nd=6�?������@ }a��?�J�LT)�?�������?5�Z(��?XV��?��Q�@�����>�?��G*�?b��Ӽ�?��jvx�?��YB���?H�z�G�?��O�V�?���;��?���˦�?Q
�C�?����1�?�G�z�?��1�2�?)�>i�??!AF��?�VYo���?������?��Q��@d��#��?����g��?�]����?P�øW�?v�=H]��?��Q���?-s��ǟ�?:�SR�?���7���??	-zռ�?��y�?�������V�o@��?�#tT��?®b�?	�e^��?�m۶m�? ףp=
�?�)�9�?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?s����`�?�0�0�?��e�s��?���]�(�?�������?ApMrx(�?}��Yc��?���_��?+��6rl�?W�m���?�G�z�	@ڨ�
�?���n��?�n0E>�?T3	Z�e�?xH����?R���Q
@�� �c�?�9vZC��?X7�"�u�?A ��X�?ƃ'��?�G�z�@��n���?�8s��?�Ox!A��?�Sq#���?/�Ij���?�G�z�@:{�N���??V�)��?_�_��?      �?��B�
�?�G�z�?�Z�K9��?��*�?9�&oe�?ߘ�[]�?��Я[[�?��(\��@%̄�?����/��?~�~��?LgR�L��?|huq���?�p=
ף�?�8G��s�?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?��Q����?�~��?O10%	s�?�M����?�G�z�׿ŝ�����?Eb���?��Y@�H�?�|��X.�?�������?��Q��	@�ڱ���?���ʦ�?�6f�@��?�~�ϓ�?FM0��>�?�G�z�@�"�T��?v��O��?��m���?G?P�e��?R��2Y��?�p=
ף@�����?)�x�?UUUUUU�?JB��EX�?�-�t�b�?q=
ףp@U��s���?~�W�f��?y@�z��?�{b�?�W�^�z�?�z�G�@�6v�KD�?b�+d�&�?�L�w�?U�&xl�?=��k�?�(\���
@?�:���?_�;I*��?k��FX�?e�5���?J����?R���Q@�A�����?���~�?9"�P9�?<O�����?!������?���(\��?�c��D��?%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�<�^�?�o��5�?O�o���?�7��ֲ�?J"���?�(\���@������?���]�?��g����?1sJJ��?��f$/��?���Q�@�T��5�?Ե7�rL�?�l��l��?���'��?��E���?��G�z��Ψ}Ri�?�v5C�?333333�?>FX�v��?$Zas ��?���Q��?�>��/��?%���y��?a8B��?�!!?�Z�?���q6�?<
ףp=�?p�n=t�?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?�
⛏A�?��P���?4 ��<�?(
P�;�?������@�X0����?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?+by,Y�?      �?B���?f���?�G�z@�1�2��?L�Q���?����S��? 0 ��?4և����?433333�?�a����?�Q���?������
@>���fi�?_*�-5�?�z�G��?� +\�?,$��?>~&.'�?      �?nt<iE��?������@�*��\�?G���;�?�x+�R�?gj��?�r4.G��?��Q�@���k>��?�>�Y��?Rb�1�?�� J`�?`�2a�?P���Q�?O|-Ϯ��?=B�k��?g�K1_h�?;9�=-�?$�D"��?q=
ףp�?�D�o��?M؜�ƹ�?x�5?,�?a�}�I<�?��Z%��?��Q��@>!R,%�?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?x����v�?4H�4H��?�)~�r��?���Kh�?�p=
ףп�����c�?����?      �?eK'b���?"�!�!��?������@��Ѐ���?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@yU�٬�?%���?G��Q
�?`�ͼ��?�Q�!\�?ףp=
�@�v#��?�&>�K��?��D/ڷ�?$�A��?�8����?֣p=
�@Q�ų5��?X���A�?������ @<�z^��?C���,�?�������?\��陌�?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?����S�?�N�u.�?�&$a��?���7�?      @6�� ��?Q�����?I�$I�$�?���Y�?z��!y�?333333�?ęmI�?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?���e��?I��/�?i�(�U�?�VC��?T���Q�?�74��q�?okL�&�?'�imt��?���
\�?۶m۶m�?��Q�@j��!��?Ŀ�y/��?.V�oD��?0�Է�N�?]2�h��?ףp=
�@�H4����?�@��+W�?��)o���?�߾���?      �?������@��&�#��?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?��]���?[�[�@�{�q�?.q����?���Q��?�@����?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�M���?��wW�?�.�E��?K^�3v�?�������?�G�z@�Z��.<�?��Lf�@�?�!��uy�?������?�aS���?�G�z@���{��?�S�����?���NV��?��=��?^���?��Q�@�D�y*��?."t��D�?]t�E�?N����Q�?�^�^�?|�G�z�?��w���?��+���?G]t�E�?X?A�x�?Ӱ�,O"�?�z�G�@����� �?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?m.���?Q^Cy�@��=,��?_�ڕ�]�?\���(\�?���^y�?T-����?UUUUUU�?L�5���?�������?ffffff @Ι�p|�?�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?#��3�U�?j|��
�?�z�G��?�����?����o.�?�(\��� @�	�x���?����,��?8�yC� @vS�+y��?K֦dmJ�?p=
ףp�6jDRf7�?�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿�_�Be�?��� ��?:��8���?��'c��?�-Wr�?333333@�)��&�?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�5�����?�������?�$I�$I@��;���?R���Q�?�z�G��?������?P@��}�?��k���?      �?�J���?�������?"t�I�+�? ��2�?S�n0�?���&�_�?I%�e��?�������?����5�?"*����?�q�q�?�s�̫~�?+1��JL�?�p=
ף�?���U�g�?/9(��?.�袋.
@�*����?�������?�������?�/%Ŷ��?������?�ol���?})3=[t�?��{a�?=
ףp=@�����?%n����?      �?7��S�?��/���?�p=
ף@�N�w��?�G,���?�	����?���R{�?��?�c��?���Q��?;⟯�:�?�r�4�?�;�;�?ڡf6�K�?�s�9��?�Q����?�+F�d��?��1���?wF]�K��?={��?������?�Q����?�K��?���,��?ى�؉��?��� W��?{�G�z�?*\���(@�)R�?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?h��Ƅ��?UUUUUU�?���t�?     ��?q=
ףp@����k��?�{㘺�?zR}%��?!�yV^�?��ծm4�?�(\���@7x�*���?��L�?��?���׈�?r�"Z�F�?���e0
�?@
ףp=�?�,>8�?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?*����Z�?48�
-�?�H�#c^�?ҞHW@�?XqBJ�e�?��(\��@��j>��?h�����?��1����?�IF��?�_{�e��?��G�zĿ� �����?���@���?��a��z�?�����?�5�3z�?H�z�G@������?�Q���?6��<�?@(��?�;�;�?أp=
�@���d�?��;��?*b�����?�0����?�8+?!��?���Q�
@���(�?��B\&�?�n0E>��?���L�?2 K��?�(\����?O(���?�l���!�?�9�s��?�1�[x}�?�[��"e�?*\���(
@�('Mh&�?�'��|-�?HT�n��?^����,�?#e�����?�(\���
@�N�8�?v��� �?o}$�o<�?��(ET��?�{i�"8�?���Q�
@��L��\�?���m,�?שǳkF�?�8��y��?@�Z���?�(\���@b��!�?-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?�X��?i�+s�?333333�?`�>��R�?��.���?q=
ףp@=�f{?��?u$_U���?7NӫT�?\:CU��?F�;�5�?433333@E����?톘��=�?+P�W
��?���gk�?�������?Z���(\�?�Q�rX��?�L���z�?X�O���?��F�{�?!���c��?�(\����?�g����?濸����?r���0�?,�C ^��?5���4�?���(\��?��ʌC�?laf"�?�q���?j�ta)��?uE]QW��?P���Q�?`P�-��?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��?������?�N��N��?��U>R
�?	f���?�G�z@�~$��?N"����?FFFFFF�?�-5��?����o�?��(\��@��2�\�?���� �?�$I�$I@W�G#��?"1ogH��?ffffff�?��a�%�?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��76�?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?^` 5��?X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?��S���?��=�9�?�[��"e�?�+U��R�?�Gq�>�?��Q���?��� g�?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿぷA�?�y�]��?]�)~I��?��@��[�?�{����?���(\�@#i��K�?dwl���?d�fI�m�?��W�6\�?=]�:��?)\���(
@^zn��?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�s����?�,B�N�?�
��v��?�߾���?������?P���Q�?z��V��?XD"���?R��+Q�?$ ����?�#F���?P���Q@]�"�H��?��B~���?ƶ#e��?-��k4�??&ǒ::�?{�G�z@8f?�?���[�?����NB�?b%c�r�?����]�?hfffff@Wd���'�?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?0�|L��?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?Ŝ�lK�?�r*��?z�Ha��?��R����?�{mĺ��?���Q�濧�7�jq�?���Y$�?��㙢�?a=]�R=�?-؂-؂�?�������?�'LZ��?�":>ɗ�?���ע�?���'-�?�R71�?      �	K�����?��H��?�z�G�?G��ֳ�?
݋н�?R���Q@X�C���?�>����?      �?0`z��Q�?'u_�?�p=
ף�?W�n��~�?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?�{Q5��?ݳ�J5��?ߣVot�?$����?�4��ǲ�?�p=
ף�?ѳ!s��?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?q�CZ�y�?)%\����??��"u��?�hJ���?433333����z��?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?�p��K"�?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?���1�^�?��;�l�?��{����?��`|��?���!�?@\���(̿Z�S�Ҳ�?(1B���?b'vb'v�?s�ӭ��? �R{���?H�z�G@K3$���?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?p;̞��?      @�њ�%g�?'u_[�?�������?y�l��?�t���?)vb'vb@nlMP��?	N�<�?�Q����?/1G��F�?n,���$�?����b)�?A�쎑��?@�1���?
ףp=
@,4�����?��Sr��?U����?<����?w�{��?<
ףp=�?�c��o�?���e(1�?      �?�KF&���?o�9)��?333333@t� �b�?B(w}1�?p�j:�?�ⷆX��?�H1�_��?���(\�@��I����?w����?     �@R���8��?�~|���?P���Q��u�%ܚ�?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?QdEc��?�����?^��?	�?�I��G�?��(\���?�~����?@i���?P��O���?�k�9���?��U�^�?(\���(�?�α	6�?����?;�;��?�(N��?�	F��?������@�ױp�9�?ۆ����?wT��~�?�f!b��?���I���?��Q�@j��+�?�4~���?h}�}-�?	+��]��?�ܽ*���?�Q���	@����P��?Sª����?      �?�	*�/�?W�<�?R���Q@[z\8s�?��_O�?��G��=�?�!|����?L��7���?033333@�P�S���?Qn�p&�?�؉�؉�?�*����?��M�`�?�p=
ף@9�>����?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�?/G�9�?�����T�?`�t����?	�m?���?��Q�@�J��}��?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?�q� .�?��"E��?�V���2�?�^�^�?�G�z�?Hݽr�?(� .b��?�k�S��?��F����?���w���? �G�z�?�&ɢ�X�?�YĘ��?9��8���?�鑢3�?^��3��?�G�z��?�*ml|��?r�2�F�?�zۜ��?z!I�,�?c[:��c�?�p=
ף@%)��a�?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�z����?��ԩ/��?AR˔���?JL �F�?�>,��?�������?���s�-�?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?M\=���?���fR�?:�:��?�Pk����?ק�����?��Q�	@WrZ~�?�����?�MA�1�?I �����?,|L���?�(\��� @����?���. �?i�`���@jڪ���?��}ylE�?�(\����?ڔ��ɣ�?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?�G����?h�[�t�?`o�3���?C�l����?
ףp=
@�T��T��?�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?��m����?�}��?       @j��_�?��¯�D�?�(\����?0-�+�?G��?�����?�8�҂�?K0�|w�?
ףp=
@�]�s��?:�"A��?��=�ĩ�?;;NL6�?���Q���?@33333ÿ�5N�m<�?|�f����?�袋.��?��q�[��?��F�?�Q���	@U5æ�)�?�.�.���?}�r��?Dw�-fV�?_�8����?8
ףp=�?���\eY�?Se�;f�?h����@A�j�}��?�WJ�B��?S���Q @���._p�?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?E� �?      �?��ԉj��?��|�nS�?333333	@��1x��?C�Z����?�Nu�w��?��سX��?�R:CW��?H�z�G@�{�͝6�?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?鄣Z��?�Dz�:�?�=��!�?���f�?�%��}'�?�p=
ף@�Ą�W�?��K_`�?      �?��]�q�?�eP*L��?R���Q@ �O���?��L��?�q�q�?G`3�!�?O���t:�?R���Q@���Bco�?����8��?��*H�?>���h�?�؊���?$\���(�?X��WI�?�O�<�?������@uq_�E�?��$2��?H�z�G�?aq8���?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?� �9�$�?h���Q��?�3�s�?�B#�E�?��Q�@� �j��?��#�N�?{�G�z�?�A+珽�?���9��?\���(\@1O�u�?R�p,C.�?������?��U�	��?n��x�>�?��Q��@���Ol�?q�ک��?      @���<X�?��=���?333333�?b�-ч�?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?It���?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?Sle�%�?Q��h��?j鱊 ��?��(C��?efffff@P�%1۶�?u��=M	�?�ڧΪu�?f>����?: 2ܫ`�?�p=
ף�?J�)f�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?�՜�pH�?�������?�m����?G��|���?E4Z����?�z�G��?hE�-\�?�j�с�?�dn}�?�xJ�Rn�?��寖�?�z�G�@�s׾�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?I��q��?�'iq��?�&��?#�����?�Q����?�E��Q�?9��%*�?�J��?N�J2�x�?*08͸�?hfffff�?���=��?�RkJ �?j��i���?��Ť��?�����?333333	@�e��O��?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?���+*�?�-шs��?���ҋ�?�#o��?q=
ףp@N�Π21�?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?��״��?Ѻ���@��O��?����T�?���(\��?���7 g�?�0�����?      @�	h�l��?t�E]t�?�p=
ף�?r��j4a�?�X$����?L�:,��?&����?G�N��?\���(�?�'�	�?���#�?��qPt�?���J��?�T�w��?�Q���?J������?
��@��?���Қ�?'::V�e�?��JR�?������	@�xE���?��TD��?x!�����?�x�;���?���&P��?�p=
ף@3�l��?�,��o*�?���tT�?Eg���?�@i�
�?��������5H<^��?���J�&�?J)��RJ�?lj�I�#�?�Y�6���?�(\���
@)����8�?�����?IM0��>�?��I��?�h�k��? R���ѿ��B+���?W['s�,�?E�JԮD�?��K�y�?��J�[��?r=
ףp@
�#�F�?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?�-J���?���|�?�o�vE��?T�P�B��?�G�z@�=�ԗ�?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?�$�l���?d!Y�B�?k���?"�?d�*|��? ףp=
׿F�w�M�?���-��?�������?�p߃���?y����?hfffff�?fd-c��?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?��ځ.��?������@GK��{��?S�<%�S�?�p=
ף�?����j��?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��?�}�!���?��Sڃ�?xE.�;	�?��}A�?��Q�@�=k,�y�?e�P���?Q`ҩy�?v����f�?2����G�?Уp=
��?6K�b0�?]��{��?�����?Iy���?E�,V!�?�Q���@�?쾕}�?�`�5^��?-iKڒ��?t��}��?Ă�� ��?�(\���
@T���%�?P��-��?�NV�#�?8��m���?�;�#�?333333@/qT��F�?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?�t&����?��(��(�?�^mSz��?g�Bg�B�?������@�5cJ�,�?��2�?�&���?YA�-��?���.�d�?�G�z@O���ii�?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�GZ<
�?�s�9��?�g�M���?���u;�?)\���(@����B�?J^��&�?���d�?���w�?�\;0��?������@3�xi��?l,����?gH���?���2G�?v�A����?�z�G��?fÿ���?�T�(Jf�?d!Y�B�?�;nRi�?��o���?=
ףp=�?��Cgm"�?S;>���?�Y���?�gS���?U�j�o�?أp=
��?���tt��?Po�S3�?!1ogH��?�8Sn�Z�?8Q�H��?�Q���@���
�S�?���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�?�k�6��?d�.���?O��N���?�UfP�h�?];0���?q=
ףp�?�⿞��?(tҶ��?�/�I��?lv��7��?��cy���?      @	���? �X��?
ףp=
�?�Ѣ�ǃ�?�;⎸#�?      @3����?�d����?���-���?_l�9��?L��N���?P���Q�?�ON���?9�KO���? ���?R-ŭX�?X�,)D�?\���(\@	`��Np�?������?v��[ʐ�?X�R5�p�?*�� 4�? �G�z���c���?��(��?7�Y�"�?ޤ�=%�?{�!���?���Q� @.�|�-0�?������?�{�D!�?�l.�VP�?�2��h.�?)\���(@���C���?��0��?R�}�=�?ӗYl�n�?.�袋.�?�Q���@N��i�?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?����?CBq�n�?�M���?ABЋf��?hfffff@?��n���?2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�V����?�SR�&�?}�K`]�?��<d��?w�C�v�?���Q�ο�*UۄP�?�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�i\|��?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�??4G0�?a�B��?�������?' Z�u�?�����?���Q�@De�&���?�]�L�b�?2&�l�?      �?]|�c���?�z�G�@h��Ơ��?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?�=�E=�?6Q�k%�?�NHL�?��{@�?T���Q�?�{�6�?�'Z�:��?�|ۗ�s�?�#%Ŀ�?�J�gQ��?��(\��@��^1���?�C����?�������?A�ra���?�@۽U��?���Q��?�/�����?���6���?�w���?zkfkl��?�k(���?      @�q�^��?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?�#jY��?z=��? ���.%�?g�#�6��?`���(\�?�w�x@�?���1�?��fy��?���N�R�?Wŵ.���?���(\�@n�-���?Jt_�h��?߈�N�@(���'<�?ZZZZZZ�?�G�z�?ۇ�����?���#�?})�Z�?d#D:��?��;�?��(\��	@���S�?�צ����?3�*�" @�#�p�j�?V�;^l	�?(\���(��9���r`�?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?�qA�[�?����=�?_r�D�Y�?�U�&�?�(\����?^ r�?�y]>d�?g;>)7�?�Ǭ�NR�?&H-/|�?=
ףp=
@VS�w �?F_L�D��?:��8���?�\�]�G�?l�����?������ @���u��?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?P�����?UUUUUU�?�k�1���?O�n�	�?��Q�@$��t�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?�C�@�?�
<h�?��+TZ�?���yV�?أp=
�@�YS����?��n �\�?�q�q�?!��s �?5/�D�)�?�p=
ף@�1Uws�?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?�_{��\�?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?�~�A
�?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?W��{3H�?mӞ��?#��~j��?�1?��l�?��i���?�Q����?Ǽ�>�?�&�j��?7��P^C�?F�����?q=
ףp�?��G�z�?:�5+�?9gήc��?�Z$�R��?������?�/��/��?033333�EF��DG�?�qV��?�z�G��?�	ϻ���?J��I���?�G�z @��w��?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�? ����?�5���?@7���$�?h/�����?�������?�y;Cb�?f�s
���?Y�%�X�?��\��?n�ٰ��? )\����?�b �*�?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?Z�yv�<�?��a�
��?��ࣹO�?:&߭��?��Q��@ ah���?O�TE���?�(፦@��x�b�?��RJ)��?�������??3�/D�?W����?��8��8�?      �?Au���?�������?(Bo*��?ݘ��2��?      �?)�gf��?B7%�!6�?��(\��տ(�~��?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?ƪ+�K�?~r!�f�?�`(vo��?l��';�?�������? !�!���?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?LG�3�K�?��=O�?M4�DM�?���2��?�ܛ���?
ףp=
@������?r+�z���?9�0s�?�~��i�?s�p5��?�G�z�@ݳ +���?����*�?)#�`��?��@�x�?�gL���?أp=
�@��ϔ��?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?:����?�5��P�?v$����?;�;��?أp=
��?�[9�.�?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?lt�&��?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff��7�z�<}�?�N"H��?����?Hx`2��?��r:���?������@�P	�_�?���q&��?      �?�ƽ7�?%Ԑ�W��?�z�G��?4�^}9�?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?!ml���?�9�n��?Ѕ�	���?��'q��?�p=
�ӿ�}G�? '�Q�^�?ᖚ�?C�7�y�?4H�4H��?���(\�@:�2�RX�?c�2��8�?l�l��?�����?T��S���?�p=
ף�? ���P��?��X��?�Kh/��?�f i5�?*g���?���Q��?{V�|4�?�מ���?�i�i�?Q�XW��?�R�~���?      �?t��3��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?Шx�?jF���?������?�.�?��?�z�G��?��2}��?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?�V��4��?]���_�?u��
	��?P�9��J�?�=
ףp�?�z�׻�?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?6%�M���?���s @N�|ҍV�?e�e��?�������?�� ��?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@��Y���?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?ű�r��?�"�hO��?���P��?��Ǹ�?���'�?�p=
ף@C���P�?9�߽9&�?(��qg	�?��K�y�?d}�OG��?���Q��?��5Pӹ�?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?QF�� �?     (�?��#qSM�?V��eЛ�?�������?�,�����?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?�����X�?t�����?�^Y�?��??��5���?ףp=
�?�!�/�?�wF�?��D'�?6������?�_�_�?�������?�Ko��?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?���@9�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?"��\��?vb'vb'�?�Mu_J�?���DxR�?���(\�ҿR��-�?+e��R�?pА����?�_P�
�?���譺�?��(\�����f��?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?�����?�NϦ�k�?�Ė��w�?���BP�?ףp=
@����?<�b���?����?�Pp���?Ŕ��%�?�p=
ף�?�����?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?��i�,�?ףp=
��?���b��?,Fڱ�?��Q�@9��V���?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�\��f��?��
�?�"nps�?�`>J�?/������?���(\�ҿ$��V�?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?t}ja>o�?\�-�=�?�Jpv��?��|j��?�������~���-�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?��F�#�?(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿�4�$��?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?���V��?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ��Ҋ��?J""}��?����;�?jZ��m�?�0�9��?��Q���?Zf����?
�&af-�??�?��?�q-���?��	�{�?أp=
��?���+��?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?W��#�^�?qCtqDbX
   n_support_qEhhK �qFh�qGRqH(KK�qIh:�C�  J   qJtqKbX
   dual_coef_qLhhK �qMh�qNRqO(KKM�qPh"�Bp  X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅���X驅����S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@�S�n@qQtqRbX
   intercept_qShhK �qTh�qURqV(KK�qWh"�C�~6~��?qXtqYbX   probA_qZhhK �q[h�q\Rq](KK�q^h"�C�:�s?�?q_tq`bX   probB_qahhK �qbh�qcRqd(KK�qeh"�C?��p@6��qftqgbX   fit_status_qhK X
   shape_fit_qiMK�qjX   _intercept_qkhhK �qlh�qmRqn(KK�qoh"�C�~6~��qptqqbX   _dual_coef_qrhhK �qsh�qtRqu(KKM�qvh"�Bp  X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?X驅���?�S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n��S�n�qwtqxbX   _sklearn_versionqyX   0.21.3qzub.