�csklearn.svm._classes
SVC
q )�q}q(X   decision_function_shapeqX   ovrqX
   break_tiesq�X   kernelqX   rbfqX   degreeqKX   gammaq	G?PbM���X   coef0q
G        X   tolqG?PbM���X   CqM�X   nuqG        X   epsilonqG        X	   shrinkingq�X   probabilityq�X
   cache_sizeqK�X   class_weightqX   balancedqX   verboseq�X   max_iterqJ����X   random_stateqK{X   _sparseq�X   n_features_in_qKX   class_weight_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�q cnumpy
dtype
q!X   f8q"K K�q#Rq$(KX   <q%NNNJ����J����K tq&b�C �?�������?q'tq(bX   classes_q)hhK �q*h�q+Rq,(KK�q-h!X   i8q.K K�q/Rq0(Kh%NNNJ����J����K tq1b�C               q2tq3bX   _gammaq4G?PbM���X   support_q5hhK �q6h�q7Rq8(KML�q9h!X   i4q:K K�q;Rq<(Kh%NNNJ����J����K tq=b�B0	              
                        !   "   #   %   &   '   (   .   /   0   2   3   6   ;   =   >   ?   @   B   E   G   H   I   J   L   O   R   X   Z   [   ^   _   c   g   h   i   j   k   l   n   s   u   v   w   x   z   ~   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �            
                          $  %  '  )  *  +  ,  1  5  9  <  =  ?  A  B  H  K  L  P  Q  S  W  X  Y  [  ]  _  a  c  d  e  h  i  j  l  p  s  u  w  y  {  |  }  ~  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                                  "  #  %  '  +  /  2  8  :  ;  @  A  C  E  F  H  I  J  K  M  O  P  S  V  W  X            F   S   V   \   o   p   {   |   �   �   �   �   �     J  ^  k    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �    !  )  -  0  B  Q  T  U  [  \  ]  ^  k  l  m  p  q  s  t  v  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                    $  %  &  '  (  )  *  +  ,  -  .  /  :  ;  =  >  ?  @  A  B  M  Q  R  S  W  a  b  c  d  e  f  g  h  i  j  k  l  m  n  o  p  q  r  s  t  u  x  y  z  {  |  }  ~    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �               q>tq?bX   support_vectors_q@hhK �qAh�qBRqC(KMLK�qDh$�B@n  �L���z�?X�O���?��F�{�?!���c��?�(\����?�g����?��=Qr�?7r#7r#�?y�sJiM�? ��c��?433333�?�Qa���?W#Q�.�?贁N�?��W9��?�$A��?!��Q��?鄣Z��?u�-BK�?��T��K�?��x���?>���~��?���Q��?f[t��?�Q���?������
@>���fi�?_*�-5�?�z�G��?� +\�?��k�<��?�k��%�?^�4�y�?��xN%�?433333�?pjh����?��״��?Ѻ���@��O��?����T�?���(\��?���7 g�?�H�^��?�i�6��?�ҩ�?���8�?Q���Q�?4�ή�5�?�5���?@7���$�?h/�����?�������?�y;Cb�?�S�����?8�P\�?��;^�?M�*g��?\���(\�?�	�;D�?�b�)U	�?�s���?�M�isT�?N1�^�?q=
ףp�?D����?�k	ԉ_�?{��z��@A�ym�?�S�r
^�?q=
ףp�?0�|L��?i�+s�?333333�?`�>��R�?��.���?q=
ףp@=�f{?��?�[{p���?�h��9�?�׻ZZ�?&*쟖1�?��(\���?��k
?�?@H�=L��?��h}�?� ��	�?Pg��)�?(\���(�??[�w(�?�j�`]�?vԥ��G�?��1_� �?��Q���?�Q����?*��Al��?4\e��?�*�z7�?a���=�?�>@,��?�z�G��?֗kx���?[��`��?ك2�*j�?� �;��?�������?�(\����?,evp��?��j�G�?u�5�o��?���d��?�~��?�G�z��?\�o�nl�?��l�
�?}+�|���?�z�6��?����6�?�p=
ף�?[�>���?���$���?�M�!�>�?�k@5�?;.l�r�?      �?�G"��?����=��?|�Zj�M�?������?���;��?�p=
ף�?��"�$��?�'=��?��fě�?��Xf[�?���¯��?�G�z @���#��?�?�}D��?��A��?!╧��?`�T�c��?H�z�G�?��1hk��?�9vZC��?X7�"�u�?A ��X�?ƃ'��?�G�z�@��n���?���\�?�^o�?�?Q�/��?^̧^̧�?�(\����?�XrYǾ�?���. �?i�`���@jڪ���?��}ylE�?�(\����?ڔ��ɣ�?��Sr��?U����?<����?w�{��?<
ףp=�?�c��o�?vP�I��?E8S8B�?������?�5��P^�?����������(�?Py�*�?333333�?@�z2;�?~r!�f�?hfffff�?�9��-c�?X��M�?      �?5T%n�?}�'}�'�?=
ףp=�?��S���?,"�j�%�?,-----�?'狗�8�?�`�����?133333�?̕x�F�?F}�p �?������?N6����?\����?ffffff�?�T����?z&�����?�H(m���?��K�y�?���cY��?��Q���?��ʦ���?��B\&�?�n0E>��?���L�?2 K��?�(\����?O(���?���RG��?"�u�)��?��s��?��o����?�z�G��?s�����?�!ފ�?c����?��J%%�?��(\���?�G�z�?�~���?f�s
���?Y�%�X�?��\��?n�ٰ��? )\����?�b �*�?/������?�k��%�?���g���?8S����?�G�z��� ���V��?�5W2V
�?<��~�?(P����?y_g6[�? ףp=
�?Q:����?��<���?      �?��(�r�?��a	G��?���(\�@n.>��	�?E�X9�x�?-��,�?)=��'�?��0���?�Q����?%ފņ,�?�O�<�?������@uq_�E�?��$2��?H�z�G�?aq8���?{J�� ��?�ǈ�d�?o���4Q�?�����? \���(�?9�IA�?�,Qʢ��?���΋��?��9�r�?�,�6
�?�z�G��?��m����?쟜�ث�?�$I�$I�?Q�d�?J��I���?0\���(�?4::RDA�?/9(��?.�袋.
@�*����?�������?�������?�/%Ŷ��?P,��v�?�������?4:�$�x�?�%����?�G�z�?Qj����?
@����?�Rǘ���?�G�y�#�?�ti'�?�Q���@c-�Gb�?{��*W��?     @�E!��p�?�$I�$��?�G�z��?�_�����?6}��a(�?)��ۘ�?*kr�/�?|�W|�W�?�G�z��?P�ϸ=�?��/����?���T4�?h�v�Q�?�����? ףp=
���A��d�?�X��S��?      �?Ѹ�U�?1�0��?���Q���rp)"���?:N�1��?G�:y�?Y<�&!�?F����?��(\���?���B�?�w�%R��?o��@�� @N�G���?�ys�%V�? ��Q��?עWG�?m��C�?      �?2zW�]6�?��L��?���(\�@��y����?Z��{��?��O ��@|cg%3�?	�<��?z�G�z�?��L�F��?$!��tN�?�+Hֹ�?:�1���?K�9���?`���(\�?K]E!�6�?�CG!�?{����D�?�/��x��?�a�a�?�p=
ף�?Щ�Y�?�%[b�F�?!t��B�?d&�X�1�?��/���?�������?y���t��?�ӄ���?R���Q@���K���?����*��?�(\����?I^J��?����o��?��p�?_�!IV�?Lx�Ie�?@
ףp=�?]T�%,u�?Ե7�rL�?�l��l��?���'��?��E���?��G�z��Ψ}Ri�?%n����?      �?7��S�?��/���?�p=
ף@�N�w��?"*����?�q�q�?�s�̫~�?+1��JL�?�p=
ף�?���U�g�?Ӡh��?a�*�Ӄ�?�{�l'K�?&c�z�u�?P���Q�?^` 5��?�S�j��?UQuUT]�?�'���?]�l��?@
ףp=�?׼����?�Պې(�?��o�j�?X�MV��?�xO�?.�?��(\���?%����?��{�A�?,˲,˲@�Z�rf�?c��0u��?���Q��?��v��?:����?�5��P�?v$����?;�;��?أp=
��?�[9�.�?(ڵ=L��?L!�i��?f��j�)�?�.6��-�?`���(\߿�4�$��?�]�`W�?J��LQ��?A���}��?��y��y�?���(\��?q0��;�?r>bܘ�?��MmjS�?e�����?|1����?���(\��?[=���?u0{UD+�?�z���?ю�hy\�?Z���/Y�?�G�z��?�ER^_1�?8����?�gS��=�?�~��H�?�Vi�_�?�������?�11�G��?���g
�?&���^B@���X^�?��FS���?G�z�G�?;��q�?z9����?#��wS	�?6��l(�?��ك	��?H�z�G�?�vף]��?�_����?      @����,��?[�o�W��?���Q��?zI%D;��? �5�0��?�����?B �Gey�?r�q��?��Q���?���I���?��;���?�`�����?��r��$�?2zh�:�?@
ףp=�?���K�?�h�(���?����?�3��=�?g�=���?�������?���w ��?_i�"�?VUUUU��?��i��?)\���(�?�������?'|im��?g�\���?�����?��񍔎�?����.��?�G�z�?'�����?�D̥�
�?�Zk����?��iz�?���\��?��Q���?��е:�?@`�ű��?����n�?sՖ$o��?h��R��?�Q����?x%�R~}�?��m��?����?&z`�5�?2u�=�S�?      �?��]�E�?l,����?gH���?���2G�?v�A����?�z�G��?fÿ���?Jt_�h��?߈�N�@(���'<�?ZZZZZZ�?�G�z�?ۇ�����?�aޤ���?�2Iw���?�ஹ��?hO�M̶�?@\���(�?���/�?&�kA�?	Q�Eΰ�?!E;q��?�������?!��Q��?��K�?L�|9��?m���X��?�B�q��?����:.�?833333�?����?."t��D�?]t�E�?N����Q�?�^�^�?|�G�z�?��w���?�
�����?���!y�?��S��?�����?������ܿ����c��?��¯e�?�Ӌ�:�?�p���?S$K��?L�z�G�?�<��2��?LH��=��?ExR��y�?���.7�?+Fڱ�?ffffff�?It���?"K�_y�?���,d�?���<�?jhɬ�?�Q���?D�&Dq�?�<�����?���Q��?��C�5�?��
=�O�?ܣp=
��?�-{X�?q����?*�3��?3iM��h�?QJ)��R�?=
ףp=�?��U#3��?��p����?      �?��e�N�?�������?R���Q@>����?���I�1�?v�ut8��?�ίZ$��?� ��^��?H�z�G�?Ґ{����?�u����?�wK�?��?�ef���?tT����?�z�G��?��-��?
�3ɦ�?�℔<��?Q澚��?�K�~���?���(\��?�`1+�H�?5-CV-I�?��;�H&�? s�_&'�?н�/B�?�z�G��?�$�(CU�?�d����?���-���?_l�9��?L��N���?P���Q�?�ON���?s����`�?�0�0�?��e�s��?���]�(�?�������?ApMrx(�?�F�,�?˕6�#��?/���K��?'i�"Ё�?�(\����?#��3�U�?J��:���?=
ףp=@��=!E�?���E�?=
ףp=�?O����?�0k��(�?�Iݗ�V�?���Y&�?���?�?      �?p��1E��?,X<`�5�?U����?D�Sj߱�?�V���*�?أp=
��?'���/��?����v
�?֤c�V��?ɰ����?���ƣ��?���Q��?ű�r��?
��Y0�?�G*;�?      �?������?��Q��?�-�����?)p�0���?2吽��?��]n�V�?�FV�a��?q=
ףp�?k^��/��?F���Ao�?�C6{ϋ�?K�Cs��?y����Q�?`���Qȿr���;�?-��#N �?����=�?j�$ŏi�?�M�4��?أp=
��?�X��?9gήc��?�Z$�R��?������?�/��/��?033333�EF��DG�?�&�j��?7��P^C�?F�����?q=
ףp�?��G�z�?:�5+�?�4��9�?��m�-��?���k���?�R~c�Q�?�(\����?�~�A
�?�[g���?B¥�K�?ñ,J�?�-�V��?أp=
��?�՜�pH�?�.YZU�?'���n"�?"�v�li�?�i��	�?ףp=
�?�X��e�?֊�q��?��Z��Z@�K��?#e�����?���Q��?
k#w��?���~���?�,�|�s�?��(��?ʁ�gA��?x=
ףp�?�k�6��?���~�?9"�P9�?<O�����?!������?���(\��?�c��D��?R�uv���?�����@�?�-�z�,�?J�a,��?P���Q�?�b�w���?�g�r�n�?|�x� �?߇�a��?�@c�Z�?@
ףp=�?�Ǔ���?�C����?�������?A�ra���?�@۽U��?���Q��?�/�����?��X��?�Kh/��?�f i5�?*g���?���Q��?{V�|4�?�מ���?�i�i�?Q�XW��?�R�~���?      �?t��3��?{��N��?""""""�?ܗ��]x�?�^Wۓ��? �G�z�?g+>����?4��Y��?���^��?	������?6���+��?|�G�z�?�<Y� Z�?�s[W��?�7�P�?Eo�h=�?�r(w��?���(\��?�TS�Yd�?�п�cX�?���؜��?��{�z��?�F��?_fffff�?�F�9���?�s���?ܶm۶m�?��xp$�?D0�i��?p�G�z�?*��g�l�?�z3��?������?{�̝{�?I�����? ףp=
�?�¹s�V�?r6]����?�������?�	��6f�?���3$��?H�z�G@��S��?*s�Z��?��r����?sڼHڃ�?�ݦz��?���Q��?-ژ���?����?u�)�Y7�?Oź1X��?9��8���?Y���(\�?���#�?��t�j�?��qg	��?d���1�?(�)��;�?�������?�O^J��?"
c���?�[�[�?��
y3�?q�M����?���Q��?�����?evoƃ��?�q�u�?�)���R�?t������?0\���(�?I��p��?�d����?��td�@�?u��s26�?�]?[��?      �?�J1�h�?�e���?R_��b#�?��L�\"�?�ԁ��0�?��Q���?A�s�я�?<�b���?����?�Pp���?Ŕ��%�?�p=
ף�?�����?0	�`���?o�vu�?N�� V�?��X���?��Q���?�/���?d��Z�?0/QzN�?g��ЯB�?㲝z��?��(\���?�}&�z�?��,���?�z�G��?����U��?a���{�?      �?KV�9d�?3�J���?�F�tj�?^���i��?�
� ��?�Q����?�\3��?���A��?w%jW�v�?Ɏ���c�?�.t���?�Q��뱿|�TT�+�?��Vc
�?x��n���?i%��G�?�oF��?�(\����?�ȣ���?D���Oz�?PuPu�?      �?٫��J�?���Q��?`d�X6�?�����?�DxR���?`f�"�?�8yh=�?q=
ףp�? ����?%˷7�	�?6�d�M6@o�辏�?ꢋ.���?�p=
ף�?�<�^�?Nɸ�o!�?���(\��?O�FG�E�?����S��?ܣp=
��?��:i�\�?/��Q��?��8��8�?�Z�_�?�������?@���Qȿg9gD�?����?k�_����?��$y���?������?��(\���?��:����?��[y��?�Ў�e��?��^*)�?z^{�?�(\����?�9)�?#
GY~�?�$�ή�?P1:BJ��?�Cc}�?q=
ףp�?�t���?����/��?~�~��?LgR�L��?|huq���?�p=
ף�?�8G��s�?9N���?�|G���?�p�Ɇ��?m��';r�?hfffff�?�p��K"�?��[�à�?��b����?��y�xi�?�cp>��?�z�G��?�)2��W�?��#���?�rcˍ-�?���'��?8��{�?@�z�G�?��'m��?K̂��?�O�պ�?�X��F�?      �?�p=
ף�?��.����?�8��;�?Ȥx�L�?h0���$�?|i�"8;�?�Q����?��H����?����� �?��(j�?�/I�a��?Dސ7��?`���Q�?��A��?�KqOq��?h�Bg�B�?�o�k��?v��/��?ףp=
�?��\���?M%����?�:�ֆi�??��!i�?��8��8�?���Q��?l�ģC�?�G��R�?�`�`�?,T����?�Cv����?���Q��?*�DXn�?��9���?�e���?��G��\�?�����\�?���(\��?:����?Un����?�������?#�R���?]�����?�Q������j;����?
�&af-�??�?��?�q-���?��	�{�?أp=
��?���+��?�,-�a��?wǋ-���?�d�?�Zց�{�?�Q����?ʞ2����?x)S�9��?�ԓ�ۥ�?!���J��?�}����?�������?������?=��*t��?�xG5���?`8����?$�Cm]�?�z�G��?��9k��?P@��}�?��k���?      �?�J���?�������?"t�I�+�?�B��w�?|�gaz�?(���t�?)��ㄍ�?��G�zĿぷA�?�?�45�?�[�[�?[�_�gx�?m�V�k�?�������?��dݔ�?��]��S�?�z�����?����?1�0��?(\���(�?j-ן�2�?������?������?�X^o�?��<t/�?H�z�G�?ȩ�*��?��2MK�?�`�`�?{���K�?�.�|��?��(\���?�٤�I��?,�,�D��?QuPu�?��a�Z�?�){�5��?���Q��?��� �?�0�1���?��8��8�?S�K�?�s����?@
ףp=�?I��~j��?fo/���?/����?'N`�4��?��3���?�������:T�+���?@�g�
�?�m۶m�@}�g?�?�%�p	�?q=
ףp�?i�o��?R8�u�?S{���?��,�1�?:�oO�$�? �G�z��S�hz���?��*�G��?t�E]t�?ؔ�
&w�?�k� ��?H�z�G�?�Gq���?0)�����?,�6z8�?�-ۗ��?�^�3=�?�������?:r����?@i���?P��O���?�k�9���?��U�^�?(\���(�?�α	6�?+e��R�?pА����?�_P�
�?���譺�?��(\�����f��?J""}��?����;�?jZ��m�?�0�9��?��Q���?Zf����?����?      �?ŵ�a��? )O��?      @�����?E�!1Y��?,1t+�?B��m��?R�(���?�G�z�?LG�3�K�?f��;��?~|`d���?|v���?�������?��G�z�?��G�A�?c&i�?�ÔP��?P>�z��?�uI�ø�?      �? ��L*r�?\�f��p�?� ���?�Z���?�Ytl�?�G�z��?[�Ӈ8�?�>H�?f�Wxe�?g��O���?&�/j�7�?�p=
ף�?�b=��
�?����?���a���?Û�P�?�`8wC�?P���Q�?���Z���?߇�WL�?~�K�`�?��,���?n�!l
�?\���(\�?�m�����?�}+>�?���?щ�z�?�2��h.�?q=
ףp�?�t�>�?U[G[��?;�;��?�	v�o�?�a�a�?������@U��A��?Шx�?jF���?������?�.�?��?�z�G��?��2}��?�(ؚ��?�{a��?Vu�o� �?      �?��(\���?T�k���?^ׅ�@�?�{a��?%�%�?yxxxxx�?t=
ףp�?�Ȳ���?�YĘ��?9��8���?�鑢3�?^��3��?�G�z��?�*ml|��?�T��?��gjƻ�?����V�?�����?\���(�?��~�qa�?szo6U��?d��֌��?8�/|p��?�Gy��?@�z�G�?���@9�?��r3��?<�A+K&�?�3i�F��?�S
�[��?أp=
��?� ;�P	�?��2���?���?��</�b�?�ռY͛�?H�z�G�?Ї�p��?�_�)���?E���K�?Mm��o��?31'��?=
ףp=�?k��f���?톘��=�?+P�W
��?���gk�?�������?Z���(\�?�Q�rX��?�fD|��?�x�3��?�Z|m��?�Hy���?@
ףp=��_��#�?c�2��8�?l�l��?�����?T��S���?�p=
ף�? ���P��?p;̞��?      @�њ�%g�?'u_[�?�������?y�l��?I@ ����?S�ѯz��?YVg�;g�?�sa�\�?(\���(�??4G0�?������?�~H���?U��oW�?��S�r
�?
ףp=
�?���y[�?1А�A�?�+��+��?+�B�i�?��	��	�?x�G�z�?<�#C��?�L�	�??q�%,�?yjBA��? k"?:��?|�G�z@�ph��?e�F-��?�������?���:%�?V���g�?ףp=
�?´�z�)�?Xe�6�?
ףp=
@�3��x�?�D�Z���?(\���(�?2�b���?�6"��t�?�[���?�r�@t �?





�?q=
ףp�?�O����?��zZ �?&jW�v%�?t���?X`��?!��Q��?���f �?��h�D��?��P��9�?�1$0��?}��O���?833333�?&~��.w�?�bf�7��?������?T���1%�?�2.ȸ�?�G�z�?�.�aq��?əPB�?��.���?gL0�h�?l��(�?ףp=
�?��m��\�?`hb&) �?'���g��?�r��o�?���%O3�?q=
ףp�?�@�I��?�_�\���?�XW.��?#�E}��?2Q覤:�?@
ףp=�?      �?�W���?{�n��?	sG�h��?в�9��?��(\���?�7���?���-��?�������?�p߃���?y����?hfffff�?fd-c��?�-��SL�?@`:�V��?��-�F�?,�~J<C�?�������?���1�^�?\	# ���?�߈��?Ľ9�X�?и[���?\���(\�?b�����?�lr����?�$I�$I�?ݗ��N�?�;⎸#�?R���Q@yU�٬�?T�.�n��?�-�׮�?H{����?������?P���Q�?��/>�?�2/۸��?�60C��? ��f��?�OZC��?�Q����?S@}�ո�?
��\���?��\AL��?)us�?      �?433333�?@�����?0�P��?��:��:�?���3f��?ѐg�:��?<
ףp=�?j��=�?5
P�j�?2ܫ`��@#'���?ߩk9���?<
ףp=�?����?O�TE���?�(፦@��x�b�?��RJ)��?�������??3�/D�?�m�02��?;r����?���	���?����<�?��(\���?�ca�M��?��{G�?����S�?Y�_��?�����B�?֣p=
��?�;S,8�?�徦�<�?�\AL� �?      �?�������?��Q��?�A���?��GA�?�6����?g�X{x�?��k(��?���Q��?=�}f-s�?�����?q=
ףp�?:D�	��?実-V��?���(\��?������?s��&�?(W�7�?���xW�?B�HV��?��(\���?�LGuk�?�𧚍��?�$I�$I@o�$���?���/��?ffffff�?9�m�.�?�1�����?UUUUUU@1��`�?n���M�?ףp=
�?�i\|��?�=>uV��?��-��-�?a#�m��?f��^�b�?D�z�G�?�V�,��?C�oB��?      �??��(b-�?b�1`�?433333@��
�f�?�M^K�?��FX��?aU]l�T�?�z8$��?W���Q�? ��Q/�?�83���?�{Nm{�?�F�� �?�������?P���Q�?1l(�?���BB�?��-b3x�?%(Ot�?ԕ��te�? )\����?��i �?�{����?�Pd����?�{c����?�������?���(\��?�ֺ��	�?6%�M���?���s @N�|ҍV�?e�e��?�������?�� ��?�!K���?)^ ���?u�`6�?���j��?q=
ףp�?(�=X��?�!ѻ�Z�?�m���V�?/�p@�p�?ve�2]��?ףp=
�?9eX��&�??d~-��?�u�����?����2�?� ?7��?      �?��Ld��?�4�i4�?,�4�rO�?�  �?���a���? ��Q��?�z����?W{�e�,�?<<<<<<�?4�,ַz�?B�:�W��?033333�?W��/.��?X���A�?������ @<�z^��?C���,�?�������?\��陌�?�h<*�?�؉�؉�?G�YH_�?�˟�Ѐ�?��Q���?��-�7�?4s���?�����?/z�V�4�?~"����?H�z�G�?��p��?��ix�?M��
���?��3�x�?���c�?x�G�z�?�0��-7�?���״�?z
!-��?���&��?\j6��b�?      �?�~�y��?O�q^�?9ÂKe�?��@�x�?*A��)�?H�z�G�?W��#�^�?5�T3�?233333@牫;X]�?�������?333333�?��W7�?��I��?      �?	)�L��?ڟ�!T�?��G�z����8I;�?�ۇA�?��*�3��?���R�]�?AA�?��(\���?���?8��?(� .b��?�k�S��?��F����?���w���? �G�z�?�&ɢ�X�?�ù�p��?+'<�ߠ�?�gdB܂�?&�}�`�?�p=
ף�?	���_�?��aJ��?��˝��?�D�y�?�$���?���(\� @��p��A�?�깘4��?�7M�?�i�'��?$p�?b�?=
ףp�\��E�%�?d�.���?O��N���?�UfP�h�?];0���?q=
ףp�?�⿞��?&1��T��?2w��!�?��WK��?t���1�?433333@�l]j� �?2�!.�?+}�G�??�sX��?�]�`#��?hfffff�?�V����?�h,�jP�?!0?N�?CޭfH��?D�#{�?!��Q��?���A��?U@�'��?�x+�R�??dM2_�?�(S�\��?�(\����B��e��?r	����?�8��8�@�m��D�?�O�?���?ףp=
��?*����Z�?aZ�/���?�p��[(�?9�����?���
b�?�������?ӆ�#�?�0�����?      @�	h�l��?t�E]t�?�p=
ף�?r��j4a�?g��5d��?�W}�p��?&I�����?�¨N���?P���Q�?�M���?A*��?�8�Mq��?E�f ��?1�C0�C�?��Q���?�M�2�?���+�? ��18�?ދ\���?I�ڸ�*�?�Q����?Rh���+�?-����?ӟ���?���;<�?�׷0���?�Q����?���e���?�,B�N�?�
��v��?�߾���?������?P���Q�?z��V��?	�F@�?�����?c�I���?l��&�l�?!��Q��?��QU��?��WJ#u�?m۶mۖ�?�t�}��?/�����?`fffff��7�z�<}�?��Ʀz��?��*�{7�?�
���?�o��o��?733333�?lt�&��?0.Ba��?.�袋.@�
�l�?haz�g�?      �?��O�^�?:+��?NB�3�?Ci!��?r�q��?Y���(\�?��F�#�?L�Q���?����S��? 0 ��?4և����?433333�?�a����?�_����?��.��@�ʌ����?�v���?��Q���?> �xka�?cL	�"��?MH�i��?'�Y&���?-K�Ӳ�?�G�z��?�Y��.�?�d�����?�T��{�?�jK?��?�"9�{�?ףp=
׿�_�Be�?8P��A��?�\;0��?<b���e�?y{�X�?      �?�`���?��V*O��?�℔<��?�vo,�q�?�쾽��?�(\����?u��׿�?��M1��?�%�8k��?�C���?�������?P���(\�?~Dk���?5~�lk��?u32"��?8����j�?�����?�z�G��?C�j���?޶z�4�?]t�E@/�_�]O�?�l�w6��?x�G�z�?g?�V.�?&�6-��?�����?d6�^3]�?��/�R/�? \���(�?D�B���?T,���?T:�g *�?"�[��t�?7.Hj��?�������?�o.�u�?*�fV=�?'���?<��v��?ZLg1���?�������?��tA���?^e�NF��?�}�K�`�?GT��a�?&Դ���?P���(\�?iS�}s��?����8��?��*H�?>���h�?�؊���?$\���(�?X��WI�?���h��?���{��?k 2-�?b�V�;��?�G�z��?9ƥ��?RWU*�?�R�?L���"��?oe�Cj��?@
ףp=�?|? ��@�?gDAl���?<e�U!�?��-��?'u_[�?�Q����?"�R[WD�?�s	��>�?��i��i@b�5:��?ܹs�Ν�?��Q���?Ŝ�lK�?�#tT��?®b�?	�e^��?�m۶m�? ףp=
�?�)�9�?�G��Q��?���|N��?#�Jc�?��� �R�?��Q��@��Y���?T�����?{NRZ��?{ʹZS��?�ϩ�~�? ףp=
ǿ��Ҋ��?��4f �?	�#����?�.�W�?]�Ib���?H
ףp=�?�	ږ@��?x�����?��S	�?NX5B���?�۷o߾�?��G�z�?W��{3H�?�.@�`�?m��;���?�kP`�^�?��u�9��?��(\���?��m e��?M�̷�?����?�Z,�0t�?8���؊�?1
ףp=�?t��Y��?�'���?�*H^�?�����?Oozӛ��?,\���(�?��x~q��?܃}����? %�2��?Z+B�߈�?�"�&o�? ףp=
�?��=�?�����?)�����?�s�H�?�u�y��?�G�z�?�!�}��?2E�Ĵ�?	��-��?'m�`�?:o1���?hfffff�?��E T�?�}�}+��??���M��?b�?O��?4CxP��? ףp=
�?կ~_�:�?�/�M�?!'n6��?U�,��#�?=��Y��??
ףp=@�s����?�_ <ʳ�?��jZǛ�?��QOy�?��paR�?      �?ӛ�L���?�t�!O�?��+��+�?��\�2�?�2����?`���(\�?�X�!)b�?�O��?v0f��#�?�3��!�?А��3$�?�(\����?vY�{4�?���6���?�w���?zkfkl��?�k(���?      @�q�^��?�WF@ �?P��^�Q�?b*d��?||9�=�?@
ףp=�?�5�����?׽�W2��?�6�i�?'�u�~�?L+0���?,\���(�?��y_���?�Ni�3�?�l�����?��+���?�S�n�?!��Q��?�{Q5��?FaAؒ�?�?<e�n�?�h�g0�?��b���?أp=
��?�_{��\�?(i�RuU�?�,˲,�@�n�*��?9��8���?���Q��?��76�?*$ȗ.�?u��GZ��?�o�k��?P��)�?�p=
ף�?���V��? Jx5��?�a�a�?�;x��<�?�������?�Q���@8)���>�?@�X兞�?f���?����15�?�>��?��Q���?r}�T��?����C��?r�Ф��?h�]8���?J�$I�$�?�G�z��?M\=���?��~���?�_��!}�?B�j
��?��XK�?      �?B9=�_��?����-�?��L��L@;K�*�O�?��
��?�������?��R{~��?�S�����?���NV��?��=��?^���?��Q�@�D�y*��?���t &�?�(��i��?����!f�?HˢBޯ�?أp=
��?�����?9�Й���?�Zs�|
�?�Ė��w�?!O	� �?�G�z��?:��]��?A��غ�?N���R�?FT~~��?�r�~��?!��Q��?����g�?�?jr~*�?       @�_ %���?��P^Cy�?�p=
ף�?�\��f��?tZQ��?I�$I�$�?�5�����?�8��8��?)\���(�?���p9�?��/f��?�^�%�?Aᚢw�?_=��Y�?:N����?J��I���?�K؞n��?Bm����?�d60Δ�?I�-U��?!5cn:�?,i�y��?ʭΛ���?ɣ��#�?x��{���?��(��?Ī����?�Lxޏ�?G�����?]fp[�	�?x5�"x�?���S(�?����>��?�������?������?7�X����?א�T�`�?�z����?�!��H'�?#<�M5��?i�(��?����#5�?f��[h��?ɗ���`�?�mKI�?8������?���D�?���Kp��?�IBb�[�?�j7���?[$g#��?@�i���?�D��N�?�V�=z� @�H�>�P�?X�b���?T" �*��?:���&�?Ӫ�Nt/�?n0���@x0��O�?�{�����?gʲ�A�?�>�����?8Z���$�?'whi.@����T�?���r���?�Î´�?A��V$�?��u��?�3��t��?
9����?����%�?^�%��.ǿ�#x�<�?C
�h�^�?y���r{�?_��֬��?p����?N����l�?�×���?�>P�!��??M��_��?7ϋ�R��?��6�x��?�@�g�M�?_!j\`�?ur��?jxAi>��?�d�A7��?�|,H�p�?#�����?�&4!S�?��Ē5��?��E�"�?z���^s�?$;(&#�?~�/1�j�?��s��?�Қ�? ��Y��?P�^���?��P��I�?}��~5��?�p���G�?w� 	��?��3K�h�?F
���f�?��L�)�?�L�y���?��Ȍl+�?0_-�?���/e�?����?�TdѮ��?����=��?�@\V�?I���� �?�c_���?�B5���?����?�D�\5��?�L44j�?z˭D}�?}bI�%�??����?�Htlݐ�?�*%SPU�?�L�G�?�r�z���?�X��z�?�nٚt�?��C���?�?�	���?I���A�?G�]�ny�?t�I	&�?�X�UA��?#��x,��?|8�:��?R4�QI�?��x����?������?.��tt�?���A�R�?����K�?�"t�b%�?,(nq���?j���2��?4�r�O��?B�㳌��?<EKE��?(�5:���?�o0V9�?]Ҵ�݀�?�\��@��?�8��y��?%)d��?�/�O�?��Ax�?��׬���?@}�)V�?��Vi�?�ĉVҎ�?�3mY��?`1����?�mG0��?��fL���?4����?��<D�?��
����?���S-��?W&+��?�\N=��?��4�<��?G
�-$��?���Ӻ�?�*^F �?��'��?⾉�=��?؝�5��?�UU�8��?��S����?�~��(�?���Y���?&������?��Bw���?F}���?�@�֑�?^��~^q�?�<e΃�?�:3��F�?�h9�m�?
�p4���?�HD��?_��Fѱ�?k�ۢd?�?�1ݪE�?}\���?IZ��?����1�?�u�)�?��_a��?��[1��?�j-e���?�Z�=��?�.�r*�?W���#�?�sP7�w�?R�[�_��?l>!�1��?ʳ�A��?!�����?ƨRZ���?��`���?�+�NNq�?y9��*��?'\���(�?MҔj�+�?E׊�ܸ�?|��XU�?�%Z�?<�<�h��?š����?��$2�?���i���?W�����?0L�rYt�?v;��D��?(\���(�?d��^a!�?����{��?}«��?�V's�?�x[9��?(\���(�?۟8t�%�?�iP��?V�����?[0�S���?�ut��z�?��]���?��<rM�?���Mۇ�?�\��?���C��?��@�?������?�n�D�-�?hi���?IJ^�^"�?�XJ)`�?��n��k�?zJ�߰��?������?:��N���?��[NE��?0@�cSQ�?t�V{F�?���5�? �9:-w�?�;Z���?��p߄X�?V�)j��?4��(���?��O0��?���)2g�?�^��?ꁣ{���?���yפ�?�2��-��?
y���?�������?��y�#�?̱G����?��B�L��?�}�p�?_�Li�0�?/лIE��?t������?�&�!��?�-�b�?+�T7�	�?��u�_��?Cl��J�?��
8|��?��X<���?��&��g�?�v`����?8A���?����C,�?d��d��?Z���K�?���R+��?��;}�?��N����?_�Y�?浲�?B:�?��DFL��?#�S���?�<�Ґ�?��0����?\Z�)��?��N���?*�x���?A�ȩ� �?&�<�0��?V|gtm
�? ��R���?�B�*�&�?%�՛��?��6���?��8��?��éa�?繛���?^"�J�G�?�\�0`��?5�p�4�?Zp:���?NA��p��?���{���?{�ov)�?����)��?�H���?؁�W�t�?U=zB�>�?�v!���?S�@�\�?���Ϊ�?B�6M�V�?&�+JΆ�?�Bp%�?�T�:���?���ST�?fh`Y#��?_�}��q�?��J=���?�L�:W�?�M���?	��	�?4I$x��?�$\xZh�?�|ߪI�?\�A?.��?�*�h/�?���vI��?�#[�?��?J��<>�?��$P��?��Bu<��?�3E�r_�?�i��X+�?Je3@�?�[+'h9�?�P^��d�?R�W}h��?_�����?��r��@�/Y{/�?�㵉��?�y��{'�?gޥ"��?��8*�Q�?� �p�@OBٺ���?Q�M�?��͓|�?p�D��9�?���)��?���G`@��K�*�?�˶�/��?�a��%�?_�3���?��|�S�?��W�@�eL]���?1U#���?�Գ���?��-U�7�?��&��?n����@\K��4�?����!�?�}kJK�?��]�4/�?�klnS�?�Nڀ�@�]Q�T��?*�cK���?j��7�?}Z4�g8�?��,�?�������?捄tk��?�"VO���?p��c���?�����d�?��]��	�?B�	�N�?d-�xi��?�:�G���?��hz9_�?��^�	�?�E<V�?H�v��?���0��?��I8���?��;�IB�?�<�*�{�?��/N��?j�����?g�)���?�8��?ӛƥ'�?G0@Rܕ�?�Q�]� �?~���D��?o7�B��?\��П�?0��9N�?B��Z�?��-0Sd�?� ��K�?�JM�VD�?�X,��?������@��t�6�?��8g�?� ��Y��?]x;�P�?����{��?��Q�\� @PDnWi�?i�5�fR�?n�����?��wִD�?��}07�?�v*�-Z @�DK�1�?��S	7u�?���3�?̦m��=�?����!l�?��#�� @����?H�<�V,�?��4�Q��?��*�o��?ڭp����?�	c��P@���C���?�r��?�eU��o�?�^�o�P�?.v����?�o���@�N/"4n�?�^7���?�d�b���?*z���V�?(9.f��?^~�!�@Uީ���?��\���?	Ip���?�I����?ֺ@"?�??�B�sſ�Kڜ+�?�dR��?*��F�_�?��-���?K'�\^�?{3�����?VJ��/�?��fR��?�ə�;��?��S����?�qKA� �?�p�Kt�?`y�0,�?�6�X��?�5��Z�?]톳K��?v�P��x�?�Wl��?�ՠQW�?��43��?�W���?2Mށ��?ˇ��E�?r,g"̥�?��e
��?���|���?�(�aU�?R!l����?Y���[�?�o���!�?9��x�H�?�ݠ{���?&�G՛�?�'�k��?�Hc�t�?m�NW�J�?��d�3��?4���9��?�M��#C�?3�����?���d�?���_���?��y[�?ƭ�����?^@��R�?FkC�{:�?���t$��?��[��?��/���?���Cv�?�γc*�?Rq(�^P�?h�� 5K�?�\�D���?
:-�<6�?��!��?�ؒ�1�?�ͫǅ5�?�۴�S��?�m\3�G�?� /��?^|�*y�?[(�P��?ڂ4	J�?S�z�+�?�o���?fm���?�D�ڴ��?��a�>�?�7�n�>�?�i~���?�4u �;�?���=T�?��	�{z�?�������?���M�?�T��j:�?Rx* *�?Db��c�?��]���?��To���?��y�4��?��)����?4oŌ�S�?���Q��?�O+���?OH����?E���b�?��!w���?�-CL@=/��f�?}ghH���?����?����?ǵ.d�j�?���jy��?Z?nS~��?e��4��?Aq#-Uo�?1AȀw�?����6W�?6m R}��?�h��6=�?�T����?R{�J��?����v�?0���9��?6P�K��?�^刦��?�a�|��?��T_E�?�_6��?Բ��[�?��wf�?��f$�?̬�f���?�>�-E��?�P�v�?���y� �?�OuD�?�����_�?�,�9�?n�˄ҁ�?�����?��R.��?tG��S�?�z&��,�?v�V�s��?�y�Wu�?
.�����?t�̥�8�?�5m���?&�c�&��?
�����?Q>}w�?2H�@/��?Zɖ���?�c�����?�.%���?�-���?�$d�ɢ�?�-�����?i��n^�?1wFB���?�y˭��?��H1���?/�{���?K��;V��?�u���'�?`��!_�?w���ѱ�?�K8s��?�秅Ч�?��R���?2��5.�?��%���?UA�bh�?t�J����?��pt@�?n����?X�	����?�J$�j��?lhƮ���?+�g�?W�����?"v5����?F�1�C�???2��?��m|0��?Y½C���?yӮj�S�?��j��t�? e8(�?m��!��?�C��8k�?Ҋ�U���?�Qq���?�L-1��?'V1�%�?p@���?-�r��?��u��?:�ș�?�����H�?}�D%0��?UԳ@�?����?K�:b��?���0�?��ä�c�?v�� ��?�՘T�?�QA�?,�K)���?1�,��?��z���?��/���?����@2�?�m}���?���H`�?�g �:��?������?F��6���?P�-���?��`?��?$�@��?o$5*|�?ϔl�@��?p��gs��?���o��?��N�o��?Ub�vC��?�/��>�?jF�#�?��7�>�?���-)��?F��X��?�K��ް�?V��"���?eȿ?�?X/�<b�?ѧf�8��?i�H�&�?K��{p'�?a�?�?�6^C�?+������?�;�����?���?�Ήx*��?q�ڄ���?y+�O	z�?_���?:��
��?4�q4�x�?������?$�ɰ'��?t�?u8`�?S
I�?��mg�?�ӗ�'T�?u����?{��>���?�l�����?/�}��?{-��B�?c���>�?��J�Hq�?�#%�-�?��'y��?������?���ڽ@%ob�G�?5���S�?��>��M�?P�¢��?"f�����?%�K��@h���]��?ѣ��M`�?.B�Z(�?�6�'�?r��%��?xP���4@�Џـf�?���z�?�{�L��?��4���?N�`a�s�?N�y�gl@��	J�$�?���`�V�?��O�ĳ�?�r`��'�?sQ���L�?�Xڪ�@��H#��?:�ƫ�?�t\JLd�?���%��?�d�
ӹ�?x$���@�fOؔ��?3�)ꦆ�?�h�c���?8�10�?@�����?��@+�N
��?n�(O�n�?%���(�?t,�	1�?��Ԡ̍�?��g@�
3���?�^��BO�?�o�Ԗ��?!U(k($�?*�6E���?@L�H\&@rwZ=��?ֈ��ו�?����?5�*��?Z?�/t��?1
f6R�?����*�?^
%���?���͋p�?^(ƩMu�?t9!1�H�?���
y�?�������?TS�w��?�	gt�?'c��?�o��W�?��sR(�?��Š���?�L+ō�?�>�7	�??��|�?wڋM��?�D5���?^��Ri;�?4�祴�?��y|ݬ�?�W�N+c�?�:ܕ"�?���cu��?sIؒGE�?jC����?Kӷ����?^��C{�?0��ne3�?�Δ�d�?��m��?@e�$���?��g�}��?͓5���?�lD4�?"0s���?dF!w��?��ˉ ��?"��b�w�?^Y-���?�(��H�?�m��8�?�P�a�Q�?��`��?Q��9�F�?Rk�J^�?~(�C�u�?��
猘�?���H�?���gm��?�x�#>N�?�g���?aV�ym1�?#��T�|�?&�ƣS�?*�n ��?�����;�?d��}��?N��'�?v���i��?���q�T�?�R�C��?=�}����?������?�/dBDe�?���?:�s$�?l)��?cO�;��?_�!p�?;	��P��?4߱E���?�����?�����:�?��j��?�a����?���	��?"���D7�?|�䛪��?�qg�\�???��+��?R;��?���̦��?�ܘ����?�܆&G�?�j4���?�����?�����?!,��_7�?����}]�?����/�?�M�89��?��Z����?ｊ�D:�?��D���?3�T���@�-l
J�?�����?�WQNc��?'j
c���?��I��?.Jy;�@�W
��??�v���?���9�??~%F���?q�Ht�?M;�&���?��H��?�_g����?(�q�\�?��s���?�hҭ�?$;;Z}@�
�%��?��R�Н�?���|���?�"���?~,�w�f�?���]��@�/}����?�n)	�?�Pg�$��?��' (��?�/��~X�?���{�f�?�z5v�?�w$� �?o��?P�?��O��?d��T�>�?3�SY);�?K��/��?!�~�-j�?b9�!1�?ˋ��Cy�?[WwwX�?w���h�?j�� �?�ׯ�=
�?�i0�f��?Թ����?�v!N��?��� �?�'�����?O��̍�?
����n�?�1���?���PS��?����]�?���B�?e0�?������?Hʮ���?�_,�P�?�:�ϱ�?[ϸ����?��}���?>�f���?� �IXn�?Qǃ<��?&\���(�?T��g&6�?Xk܃�?��H��t�?����%��?N��;Ru�?!��Q��?��W��;�?ܳ��"�?�@Gn��?*x�dv��?�����?�����? ���j2�?�s���?�������?Ԅ�����?w߅>��?�+7���?S��8\�?E����?��nT��?��
0��?Ә�H5t�?�96=��?����1�?vs�ɗ��?';���?��$��x�?��c�}_�?Q�7��?�L���
�?.
U�?�?#��~9@��,��V�?7�EҚ��?[E-yY�?�����?�τ�!�?qR�nQ�?1d�{��?e��O��?�pW8'�?8
��j�?��y���?K�$��?�?3�5<L��?#MEl��?'ñ�7�?8U ���?��g؍�?})t���?K����P�?��=p�?A�5}�?� ����?Ł#Ƶ�?���:��?=@�����?z�
� s�?30Z���?H`�'�?�3�3(�?5c0ɽ��?8�
���?���Z��?ܞ8�n�?O��6	�?�ad&��?�}�\���?mz!Ġ�?�
����?/#�v��?�`?��#�?�Ş���?9qc����?cS�q��?,�+B���?ۺ%N�?gnbg�?�ۿZ��?��.:I�?�`^P�? i՚n�?��kWr�?�Y,�E��?�r�i��?B��A�?{�v7���?l72ý�?�W��B=�?��~�8��?Am��/F�?�K���@Q�DI�?;�Lr���?}}����?/&��͡�?���W�C�?����t�@�[�5���?\=��.��?Eh  </�?�K��u�?�é���?yrn�*`@7w�@�?�;�hu�?d�.~��?M�G��(�?S��>T�?R��`��@kH��?04h��?���aH��?��m��?�3w�e��?�3QP@�|�<�B�?��J�M�?�V)	��?�\����?�����?j���y@��h���?(�=��?D�T��?��Q�OB�?(~_\C�?X�W��@���Y�?�y����?�ZQ��?��G�V�?e{��"�?k1&M���?�r�Z��?��T����?�|oKD/�?��>jl�?w&��	�?��7�N��?m7tt,��?�<?S�J�?1cE���?��
��?�k�Y��?'�l�O�?���EL�?"(ͫ�6�?���}� �?��m��c�?Ш��_*�?�j�#��?M���դ�?Lja`���?Cyit[�?�ax:R�?��}�?҅L`��?>d����?, �E�=�?��o�/��?t�"�T�?n�R�-�?��Ǵ��?�����?����7.�?�ną��?K~�߈{�?�n1OW'�?�@�x���?��}fɥ�?S�>��/�?�� y�H�?ڟ����?������?�{#����?H57O��?=�s���?��ϣ�?nM:/@�??�o)�?��_K���?���X��?.KI��?��}�?z:23f�?�nt�ģ�?���M�?�Ѳ����?ZHS�J�? d,��@���N�@�?��I��+�?0*	T�?$��һN�?�ߴ���?4����@Z�EU���?p����c�?=O\���?���7�,�?�����?���l@J��L�<�?��V��?N��S�J�?u�N�?bk$����?a���w=@?nT}���?QG1R���?���,�h�?��W��&�?6ܿ<���?�ܱ�`�@v.#~ę�?'�58�5�?l��(n��?�?;��J�?�kN�h�?���(�� @W55�6M�?��3���?q�u^�h�?v.�ܦ�?�Zma&�?�\P~��?��D����?_�|�4d�?b�D�7�?�:"�(�?���_��?D�(Ad�@�JG\���?��I��?��m�aF�?�����?�g���?i�p�L��?�6���`�?��<����?iR"����?�e����?{�����?��3�2�?�+���?.3�W{s�?��ta�?�Q?@R�?���IV�?�z�=��?�(]o&�?�?<_v�?޴D�H(�?���LP�?!��J�??� ��?���c7�?�Z3j� �?�Wg��v�?�?:����?�8�����?�S�2�?�_?x�H�?rԄ�}�?���9���?CT�X �?m?�O���?~q�'���?4(>1�?h݅6��?%hV�C�?�}�\��?�n���?�I��D^�?mjg 2��?���� �?1�aJ���?\������?�~�	"�?/��EJ�?����/Y�?���6��?�� B��?������?��G�L�?3j�.�*�?f��M`�?��Lw�
�?��έ�?�\=#��?�����I�?ym�36��?*��lF��?_�9��?��%�r��?��g���?�o�����?���E�?=sR��&�?�6|��?�h?x�w�?�b:9��?k��:�?�i��a�?cŏ �4�?(6SZ9�?�c;����?��Z��?�]uq��?��!��o�?��'���?�¨�&�?����N�?�%�G��?��Q�?��?V^8��h�?��\ݥ�?��!+��?���3+�?�;_���?�����?�� F�V�?�+��k��?U�)�С�?^�N���?S�K�&�?�~���f�?��?�w<����?ʩ�V�?]^h"�n�?�.�'��?0�O4�?�?���>��?4��'��?��$EZ�?^�d	���?� 	!���? ���?O�k����?��o�d�?������?��%� @M��X��?�#��K�?��Ѭ�?��ɷ*x�?�/�#�9�?E몆�.@UE�	��?�R�cr��?-1pM��?\u�w�i�?����0�?t�8ٜ�@��
�zO�?yo��D��?w� ���?�쬠�8�?�{ڏ��?L�ώ�@�~bh�?�6	ĜV�?��޾nr�?��:��?׭�����? �~���@	GW}<�?���8��?`̠��?݈r���?/I|���?L�-��?�?��X�L�?�N]����?Ζ���?������?��~q���?�F)�H@k�f���?�K�(�W�?�����?���b �?q(6�+��?���W(��??�t'��?trЧk�? }�\8K@q������?*�|y���?1.s��?����v��?�J����?����u@���X���?���UC�?��f�F��?#���d�?���:�?{츓@Y��U_�?G�E\g��?�D���?D�_G�Z�?���'l�?P�寠�@3�����?F�r�D��?<1c�m�?������?JV<S�?��y��� @���?����?(�x�1 @������?/���	�?���1o:�?�%^�t��?q�����?���� @�Φu[��?R`�2c�?oܯWT�?M��F ��?��t�4�?��6���?P	�>e�?� n��?��t���?����_�? �]Ro5�?x���@y��b��?JB[j��?�2�ů��?�gS#8�?LL�P� �?�J�K�@��m�1-�?����?xUz[:_�?x[`�2�?��Z<d�?,u�TX�@�>|N�O�?�"}hBp�?��p#c��?"pۘ��?8��-�?��2Hr�@r���v#�?W��?��?���Q�L�?�vI�(�? �6B��?f���?@@ȏT2�O�?l��s>�?b ���C�?Ȝ�s:�?S�F����?�Zd���?}����?��$����?�d_\�o�?���-��?�0����?2�-*�?�k�aP�?���Ca�?�_��H
�?�݇/R�?��<���?Wmʫ��?XG�D�v�?_�G+��? ���J��?6Ǚk���?�F����?i�����?���(M�?�S���{�?W�}~�z�?C�9�?�������?�Y["<�?��	y�?ݝ�ʉ�?2M��q�?M�Wو�?7����?��pT�?]z�{�?�������?�8�7���?�~����?�Y����?n�>i�?>!᧲��?Fa}�0�?R�m�%��?����z�?�&׵�)�?��u�F��?�â@�?��#Q\��?�8��q��?���V���?6�4�U�?��_{� @������?��2B��?�W�jG�?8���m�?�3_ �?5��at��?M��v`��?�a�.��?G�)�?R�q̧��?� +[�?�ұ� �?������?�����?&\���h�?�W���I�?P���	�?�&2��?��1���?��~XԢ�?Vl'<�?����61�?�� N�?�kYd�� @�ө̯�?	ܰrv�?�������?Q^a��?w!�_��?$�ѡ��?��7&�?�a��1��?�'����?�9�?Ɉ�����?c~���]�?�p�w�5�?������?��5E�R�?������?��ӛ�?;�w� @6ݩ+#m�?!���t�?∨�u��?������?�1!�_J�?e^�v�|�?&u�g��?�{B����?��B�_��?�u:�2��?�j/��s�?�tYK�Q�?�� ށ�?gFi���?L�����?��}\*�?qEtqFbX
   _n_supportqGhhK �qHh�qIRqJ(KK�qKh<�C$  (  qLtqMbX
   dual_coef_qNhhK �qOh�qPRqQ(KKML�qRh$�B`  �ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~����M�[_��ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~��������ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~��/�\�BG��ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~���ӧO�~������W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@^�--yh@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@�)oxMd@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@����W�@qStqTbX
   intercept_qUhhK �qVh�qWRqX(KK�qYh$�C��>.j 1�qZtq[bX   _probAq\hhK �q]h�q^Rq_(KK�q`h$�CDh`��F�qatqbbX   _probBqchhK �qdh�qeRqf(KK�qgh$�Co��$#+��qhtqibX   fit_status_qjK X
   shape_fit_qkMK�qlX   _intercept_qmhhK �qnh�qoRqp(KK�qqh$�C��>.j 1@qrtqsbX   _dual_coef_qthhK �quh�qvRqw(KKML�qxh$�B`  �ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@��M�[_@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@����@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@/�\�BG@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@�ӧO�~�@����W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W��^�--yh�����W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W���)oxMd�����W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W������W��qytqzbX   _sklearn_versionq{X   0.23.1q|ub.